library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;



entity rom_non_linear_mapper is
port ( 
	i_clk : in std_logic;
	i_addr : in std_logic_vector(11 downto 0);
	o_data : out std_logic_vector(11 downto 0)
);
end rom_non_linear_mapper;

architecture Behavioral of rom_non_linear_mapper is

TYPE ARRAY_ROM is array (natural range<>) of std_logic_vector(11 downto 0);

signal rom_data :ARRAY_ROM(4095 downto 0);

attribute RAM_STYLE : string;
attribute RAM_STYLE of rom_data: signal is "BLOCK";

begin


rom_data(0) <= "000000000000";
rom_data(1) <= "000000000000";
rom_data(2) <= "000000000000";
rom_data(3) <= "000000000000";
rom_data(4) <= "000000000000";
rom_data(5) <= "000000000000";
rom_data(6) <= "000000000000";
rom_data(7) <= "000000000000";
rom_data(8) <= "000000000000";
rom_data(9) <= "000000000000";
rom_data(10) <= "000000000000";
rom_data(11) <= "000000000000";
rom_data(12) <= "000000000000";
rom_data(13) <= "000000000000";
rom_data(14) <= "000000000000";
rom_data(15) <= "000000000000";
rom_data(16) <= "000000000000";
rom_data(17) <= "000000000000";
rom_data(18) <= "000000000000";
rom_data(19) <= "000000000000";
rom_data(20) <= "000000000000";
rom_data(21) <= "000000000000";
rom_data(22) <= "000000000000";
rom_data(23) <= "000000000000";
rom_data(24) <= "000000000000";
rom_data(25) <= "000000000000";
rom_data(26) <= "000000000000";
rom_data(27) <= "000000000000";
rom_data(28) <= "000000000000";
rom_data(29) <= "000000000000";
rom_data(30) <= "000000000000";
rom_data(31) <= "000000000000";
rom_data(32) <= "000000000000";
rom_data(33) <= "000000000000";
rom_data(34) <= "000000000000";
rom_data(35) <= "000000000000";
rom_data(36) <= "000000000000";
rom_data(37) <= "000000000000";
rom_data(38) <= "000000000000";
rom_data(39) <= "000000000000";
rom_data(40) <= "000000000000";
rom_data(41) <= "000000000000";
rom_data(42) <= "000000000000";
rom_data(43) <= "000000000000";
rom_data(44) <= "000000000000";
rom_data(45) <= "000000000000";
rom_data(46) <= "000000000000";
rom_data(47) <= "000000000000";
rom_data(48) <= "000000000000";
rom_data(49) <= "000000000000";
rom_data(50) <= "000000000000";
rom_data(51) <= "000000000000";
rom_data(52) <= "000000000000";
rom_data(53) <= "000000000000";
rom_data(54) <= "000000000000";
rom_data(55) <= "000000000000";
rom_data(56) <= "000000000000";
rom_data(57) <= "000000000000";
rom_data(58) <= "000000000000";
rom_data(59) <= "000000000000";
rom_data(60) <= "000000000000";
rom_data(61) <= "000000000000";
rom_data(62) <= "000000000000";
rom_data(63) <= "000000000000";
rom_data(64) <= "000000000001";
rom_data(65) <= "000000000001";
rom_data(66) <= "000000000001";
rom_data(67) <= "000000000001";
rom_data(68) <= "000000000001";
rom_data(69) <= "000000000001";
rom_data(70) <= "000000000001";
rom_data(71) <= "000000000001";
rom_data(72) <= "000000000001";
rom_data(73) <= "000000000001";
rom_data(74) <= "000000000001";
rom_data(75) <= "000000000001";
rom_data(76) <= "000000000001";
rom_data(77) <= "000000000001";
rom_data(78) <= "000000000001";
rom_data(79) <= "000000000001";
rom_data(80) <= "000000000001";
rom_data(81) <= "000000000001";
rom_data(82) <= "000000000001";
rom_data(83) <= "000000000001";
rom_data(84) <= "000000000001";
rom_data(85) <= "000000000001";
rom_data(86) <= "000000000001";
rom_data(87) <= "000000000001";
rom_data(88) <= "000000000001";
rom_data(89) <= "000000000001";
rom_data(90) <= "000000000001";
rom_data(91) <= "000000000010";
rom_data(92) <= "000000000010";
rom_data(93) <= "000000000010";
rom_data(94) <= "000000000010";
rom_data(95) <= "000000000010";
rom_data(96) <= "000000000010";
rom_data(97) <= "000000000010";
rom_data(98) <= "000000000010";
rom_data(99) <= "000000000010";
rom_data(100) <= "000000000010";
rom_data(101) <= "000000000010";
rom_data(102) <= "000000000010";
rom_data(103) <= "000000000010";
rom_data(104) <= "000000000010";
rom_data(105) <= "000000000010";
rom_data(106) <= "000000000010";
rom_data(107) <= "000000000010";
rom_data(108) <= "000000000010";
rom_data(109) <= "000000000010";
rom_data(110) <= "000000000010";
rom_data(111) <= "000000000011";
rom_data(112) <= "000000000011";
rom_data(113) <= "000000000011";
rom_data(114) <= "000000000011";
rom_data(115) <= "000000000011";
rom_data(116) <= "000000000011";
rom_data(117) <= "000000000011";
rom_data(118) <= "000000000011";
rom_data(119) <= "000000000011";
rom_data(120) <= "000000000011";
rom_data(121) <= "000000000011";
rom_data(122) <= "000000000011";
rom_data(123) <= "000000000011";
rom_data(124) <= "000000000011";
rom_data(125) <= "000000000011";
rom_data(126) <= "000000000011";
rom_data(127) <= "000000000011";
rom_data(128) <= "000000000100";
rom_data(129) <= "000000000100";
rom_data(130) <= "000000000100";
rom_data(131) <= "000000000100";
rom_data(132) <= "000000000100";
rom_data(133) <= "000000000100";
rom_data(134) <= "000000000100";
rom_data(135) <= "000000000100";
rom_data(136) <= "000000000100";
rom_data(137) <= "000000000100";
rom_data(138) <= "000000000100";
rom_data(139) <= "000000000100";
rom_data(140) <= "000000000100";
rom_data(141) <= "000000000100";
rom_data(142) <= "000000000100";
rom_data(143) <= "000000000100";
rom_data(144) <= "000000000101";
rom_data(145) <= "000000000101";
rom_data(146) <= "000000000101";
rom_data(147) <= "000000000101";
rom_data(148) <= "000000000101";
rom_data(149) <= "000000000101";
rom_data(150) <= "000000000101";
rom_data(151) <= "000000000101";
rom_data(152) <= "000000000101";
rom_data(153) <= "000000000101";
rom_data(154) <= "000000000101";
rom_data(155) <= "000000000101";
rom_data(156) <= "000000000101";
rom_data(157) <= "000000000110";
rom_data(158) <= "000000000110";
rom_data(159) <= "000000000110";
rom_data(160) <= "000000000110";
rom_data(161) <= "000000000110";
rom_data(162) <= "000000000110";
rom_data(163) <= "000000000110";
rom_data(164) <= "000000000110";
rom_data(165) <= "000000000110";
rom_data(166) <= "000000000110";
rom_data(167) <= "000000000110";
rom_data(168) <= "000000000110";
rom_data(169) <= "000000000110";
rom_data(170) <= "000000000111";
rom_data(171) <= "000000000111";
rom_data(172) <= "000000000111";
rom_data(173) <= "000000000111";
rom_data(174) <= "000000000111";
rom_data(175) <= "000000000111";
rom_data(176) <= "000000000111";
rom_data(177) <= "000000000111";
rom_data(178) <= "000000000111";
rom_data(179) <= "000000000111";
rom_data(180) <= "000000000111";
rom_data(181) <= "000000001000";
rom_data(182) <= "000000001000";
rom_data(183) <= "000000001000";
rom_data(184) <= "000000001000";
rom_data(185) <= "000000001000";
rom_data(186) <= "000000001000";
rom_data(187) <= "000000001000";
rom_data(188) <= "000000001000";
rom_data(189) <= "000000001000";
rom_data(190) <= "000000001000";
rom_data(191) <= "000000001000";
rom_data(192) <= "000000001001";
rom_data(193) <= "000000001001";
rom_data(194) <= "000000001001";
rom_data(195) <= "000000001001";
rom_data(196) <= "000000001001";
rom_data(197) <= "000000001001";
rom_data(198) <= "000000001001";
rom_data(199) <= "000000001001";
rom_data(200) <= "000000001001";
rom_data(201) <= "000000001001";
rom_data(202) <= "000000001001";
rom_data(203) <= "000000001010";
rom_data(204) <= "000000001010";
rom_data(205) <= "000000001010";
rom_data(206) <= "000000001010";
rom_data(207) <= "000000001010";
rom_data(208) <= "000000001010";
rom_data(209) <= "000000001010";
rom_data(210) <= "000000001010";
rom_data(211) <= "000000001010";
rom_data(212) <= "000000001010";
rom_data(213) <= "000000001011";
rom_data(214) <= "000000001011";
rom_data(215) <= "000000001011";
rom_data(216) <= "000000001011";
rom_data(217) <= "000000001011";
rom_data(218) <= "000000001011";
rom_data(219) <= "000000001011";
rom_data(220) <= "000000001011";
rom_data(221) <= "000000001011";
rom_data(222) <= "000000001100";
rom_data(223) <= "000000001100";
rom_data(224) <= "000000001100";
rom_data(225) <= "000000001100";
rom_data(226) <= "000000001100";
rom_data(227) <= "000000001100";
rom_data(228) <= "000000001100";
rom_data(229) <= "000000001100";
rom_data(230) <= "000000001100";
rom_data(231) <= "000000001101";
rom_data(232) <= "000000001101";
rom_data(233) <= "000000001101";
rom_data(234) <= "000000001101";
rom_data(235) <= "000000001101";
rom_data(236) <= "000000001101";
rom_data(237) <= "000000001101";
rom_data(238) <= "000000001101";
rom_data(239) <= "000000001101";
rom_data(240) <= "000000001110";
rom_data(241) <= "000000001110";
rom_data(242) <= "000000001110";
rom_data(243) <= "000000001110";
rom_data(244) <= "000000001110";
rom_data(245) <= "000000001110";
rom_data(246) <= "000000001110";
rom_data(247) <= "000000001110";
rom_data(248) <= "000000001111";
rom_data(249) <= "000000001111";
rom_data(250) <= "000000001111";
rom_data(251) <= "000000001111";
rom_data(252) <= "000000001111";
rom_data(253) <= "000000001111";
rom_data(254) <= "000000001111";
rom_data(255) <= "000000001111";
rom_data(256) <= "000000010000";
rom_data(257) <= "000000010000";
rom_data(258) <= "000000010000";
rom_data(259) <= "000000010000";
rom_data(260) <= "000000010000";
rom_data(261) <= "000000010000";
rom_data(262) <= "000000010000";
rom_data(263) <= "000000010000";
rom_data(264) <= "000000010001";
rom_data(265) <= "000000010001";
rom_data(266) <= "000000010001";
rom_data(267) <= "000000010001";
rom_data(268) <= "000000010001";
rom_data(269) <= "000000010001";
rom_data(270) <= "000000010001";
rom_data(271) <= "000000010001";
rom_data(272) <= "000000010010";
rom_data(273) <= "000000010010";
rom_data(274) <= "000000010010";
rom_data(275) <= "000000010010";
rom_data(276) <= "000000010010";
rom_data(277) <= "000000010010";
rom_data(278) <= "000000010010";
rom_data(279) <= "000000010011";
rom_data(280) <= "000000010011";
rom_data(281) <= "000000010011";
rom_data(282) <= "000000010011";
rom_data(283) <= "000000010011";
rom_data(284) <= "000000010011";
rom_data(285) <= "000000010011";
rom_data(286) <= "000000010011";
rom_data(287) <= "000000010100";
rom_data(288) <= "000000010100";
rom_data(289) <= "000000010100";
rom_data(290) <= "000000010100";
rom_data(291) <= "000000010100";
rom_data(292) <= "000000010100";
rom_data(293) <= "000000010100";
rom_data(294) <= "000000010101";
rom_data(295) <= "000000010101";
rom_data(296) <= "000000010101";
rom_data(297) <= "000000010101";
rom_data(298) <= "000000010101";
rom_data(299) <= "000000010101";
rom_data(300) <= "000000010101";
rom_data(301) <= "000000010110";
rom_data(302) <= "000000010110";
rom_data(303) <= "000000010110";
rom_data(304) <= "000000010110";
rom_data(305) <= "000000010110";
rom_data(306) <= "000000010110";
rom_data(307) <= "000000010111";
rom_data(308) <= "000000010111";
rom_data(309) <= "000000010111";
rom_data(310) <= "000000010111";
rom_data(311) <= "000000010111";
rom_data(312) <= "000000010111";
rom_data(313) <= "000000010111";
rom_data(314) <= "000000011000";
rom_data(315) <= "000000011000";
rom_data(316) <= "000000011000";
rom_data(317) <= "000000011000";
rom_data(318) <= "000000011000";
rom_data(319) <= "000000011000";
rom_data(320) <= "000000011001";
rom_data(321) <= "000000011001";
rom_data(322) <= "000000011001";
rom_data(323) <= "000000011001";
rom_data(324) <= "000000011001";
rom_data(325) <= "000000011001";
rom_data(326) <= "000000011001";
rom_data(327) <= "000000011010";
rom_data(328) <= "000000011010";
rom_data(329) <= "000000011010";
rom_data(330) <= "000000011010";
rom_data(331) <= "000000011010";
rom_data(332) <= "000000011010";
rom_data(333) <= "000000011011";
rom_data(334) <= "000000011011";
rom_data(335) <= "000000011011";
rom_data(336) <= "000000011011";
rom_data(337) <= "000000011011";
rom_data(338) <= "000000011011";
rom_data(339) <= "000000011100";
rom_data(340) <= "000000011100";
rom_data(341) <= "000000011100";
rom_data(342) <= "000000011100";
rom_data(343) <= "000000011100";
rom_data(344) <= "000000011100";
rom_data(345) <= "000000011101";
rom_data(346) <= "000000011101";
rom_data(347) <= "000000011101";
rom_data(348) <= "000000011101";
rom_data(349) <= "000000011101";
rom_data(350) <= "000000011101";
rom_data(351) <= "000000011110";
rom_data(352) <= "000000011110";
rom_data(353) <= "000000011110";
rom_data(354) <= "000000011110";
rom_data(355) <= "000000011110";
rom_data(356) <= "000000011110";
rom_data(357) <= "000000011111";
rom_data(358) <= "000000011111";
rom_data(359) <= "000000011111";
rom_data(360) <= "000000011111";
rom_data(361) <= "000000011111";
rom_data(362) <= "000000100000";
rom_data(363) <= "000000100000";
rom_data(364) <= "000000100000";
rom_data(365) <= "000000100000";
rom_data(366) <= "000000100000";
rom_data(367) <= "000000100000";
rom_data(368) <= "000000100001";
rom_data(369) <= "000000100001";
rom_data(370) <= "000000100001";
rom_data(371) <= "000000100001";
rom_data(372) <= "000000100001";
rom_data(373) <= "000000100001";
rom_data(374) <= "000000100010";
rom_data(375) <= "000000100010";
rom_data(376) <= "000000100010";
rom_data(377) <= "000000100010";
rom_data(378) <= "000000100010";
rom_data(379) <= "000000100011";
rom_data(380) <= "000000100011";
rom_data(381) <= "000000100011";
rom_data(382) <= "000000100011";
rom_data(383) <= "000000100011";
rom_data(384) <= "000000100100";
rom_data(385) <= "000000100100";
rom_data(386) <= "000000100100";
rom_data(387) <= "000000100100";
rom_data(388) <= "000000100100";
rom_data(389) <= "000000100100";
rom_data(390) <= "000000100101";
rom_data(391) <= "000000100101";
rom_data(392) <= "000000100101";
rom_data(393) <= "000000100101";
rom_data(394) <= "000000100101";
rom_data(395) <= "000000100110";
rom_data(396) <= "000000100110";
rom_data(397) <= "000000100110";
rom_data(398) <= "000000100110";
rom_data(399) <= "000000100110";
rom_data(400) <= "000000100111";
rom_data(401) <= "000000100111";
rom_data(402) <= "000000100111";
rom_data(403) <= "000000100111";
rom_data(404) <= "000000100111";
rom_data(405) <= "000000101000";
rom_data(406) <= "000000101000";
rom_data(407) <= "000000101000";
rom_data(408) <= "000000101000";
rom_data(409) <= "000000101000";
rom_data(410) <= "000000101001";
rom_data(411) <= "000000101001";
rom_data(412) <= "000000101001";
rom_data(413) <= "000000101001";
rom_data(414) <= "000000101001";
rom_data(415) <= "000000101010";
rom_data(416) <= "000000101010";
rom_data(417) <= "000000101010";
rom_data(418) <= "000000101010";
rom_data(419) <= "000000101010";
rom_data(420) <= "000000101011";
rom_data(421) <= "000000101011";
rom_data(422) <= "000000101011";
rom_data(423) <= "000000101011";
rom_data(424) <= "000000101011";
rom_data(425) <= "000000101100";
rom_data(426) <= "000000101100";
rom_data(427) <= "000000101100";
rom_data(428) <= "000000101100";
rom_data(429) <= "000000101100";
rom_data(430) <= "000000101101";
rom_data(431) <= "000000101101";
rom_data(432) <= "000000101101";
rom_data(433) <= "000000101101";
rom_data(434) <= "000000101101";
rom_data(435) <= "000000101110";
rom_data(436) <= "000000101110";
rom_data(437) <= "000000101110";
rom_data(438) <= "000000101110";
rom_data(439) <= "000000101111";
rom_data(440) <= "000000101111";
rom_data(441) <= "000000101111";
rom_data(442) <= "000000101111";
rom_data(443) <= "000000101111";
rom_data(444) <= "000000110000";
rom_data(445) <= "000000110000";
rom_data(446) <= "000000110000";
rom_data(447) <= "000000110000";
rom_data(448) <= "000000110001";
rom_data(449) <= "000000110001";
rom_data(450) <= "000000110001";
rom_data(451) <= "000000110001";
rom_data(452) <= "000000110001";
rom_data(453) <= "000000110010";
rom_data(454) <= "000000110010";
rom_data(455) <= "000000110010";
rom_data(456) <= "000000110010";
rom_data(457) <= "000000110011";
rom_data(458) <= "000000110011";
rom_data(459) <= "000000110011";
rom_data(460) <= "000000110011";
rom_data(461) <= "000000110011";
rom_data(462) <= "000000110100";
rom_data(463) <= "000000110100";
rom_data(464) <= "000000110100";
rom_data(465) <= "000000110100";
rom_data(466) <= "000000110101";
rom_data(467) <= "000000110101";
rom_data(468) <= "000000110101";
rom_data(469) <= "000000110101";
rom_data(470) <= "000000110101";
rom_data(471) <= "000000110110";
rom_data(472) <= "000000110110";
rom_data(473) <= "000000110110";
rom_data(474) <= "000000110110";
rom_data(475) <= "000000110111";
rom_data(476) <= "000000110111";
rom_data(477) <= "000000110111";
rom_data(478) <= "000000110111";
rom_data(479) <= "000000111000";
rom_data(480) <= "000000111000";
rom_data(481) <= "000000111000";
rom_data(482) <= "000000111000";
rom_data(483) <= "000000111000";
rom_data(484) <= "000000111001";
rom_data(485) <= "000000111001";
rom_data(486) <= "000000111001";
rom_data(487) <= "000000111001";
rom_data(488) <= "000000111010";
rom_data(489) <= "000000111010";
rom_data(490) <= "000000111010";
rom_data(491) <= "000000111010";
rom_data(492) <= "000000111011";
rom_data(493) <= "000000111011";
rom_data(494) <= "000000111011";
rom_data(495) <= "000000111011";
rom_data(496) <= "000000111100";
rom_data(497) <= "000000111100";
rom_data(498) <= "000000111100";
rom_data(499) <= "000000111100";
rom_data(500) <= "000000111101";
rom_data(501) <= "000000111101";
rom_data(502) <= "000000111101";
rom_data(503) <= "000000111101";
rom_data(504) <= "000000111110";
rom_data(505) <= "000000111110";
rom_data(506) <= "000000111110";
rom_data(507) <= "000000111110";
rom_data(508) <= "000000111111";
rom_data(509) <= "000000111111";
rom_data(510) <= "000000111111";
rom_data(511) <= "000000111111";
rom_data(512) <= "000001000000";
rom_data(513) <= "000001000000";
rom_data(514) <= "000001000000";
rom_data(515) <= "000001000000";
rom_data(516) <= "000001000001";
rom_data(517) <= "000001000001";
rom_data(518) <= "000001000001";
rom_data(519) <= "000001000001";
rom_data(520) <= "000001000010";
rom_data(521) <= "000001000010";
rom_data(522) <= "000001000010";
rom_data(523) <= "000001000010";
rom_data(524) <= "000001000011";
rom_data(525) <= "000001000011";
rom_data(526) <= "000001000011";
rom_data(527) <= "000001000011";
rom_data(528) <= "000001000100";
rom_data(529) <= "000001000100";
rom_data(530) <= "000001000100";
rom_data(531) <= "000001000100";
rom_data(532) <= "000001000101";
rom_data(533) <= "000001000101";
rom_data(534) <= "000001000101";
rom_data(535) <= "000001000101";
rom_data(536) <= "000001000110";
rom_data(537) <= "000001000110";
rom_data(538) <= "000001000110";
rom_data(539) <= "000001000110";
rom_data(540) <= "000001000111";
rom_data(541) <= "000001000111";
rom_data(542) <= "000001000111";
rom_data(543) <= "000001001000";
rom_data(544) <= "000001001000";
rom_data(545) <= "000001001000";
rom_data(546) <= "000001001000";
rom_data(547) <= "000001001001";
rom_data(548) <= "000001001001";
rom_data(549) <= "000001001001";
rom_data(550) <= "000001001001";
rom_data(551) <= "000001001010";
rom_data(552) <= "000001001010";
rom_data(553) <= "000001001010";
rom_data(554) <= "000001001010";
rom_data(555) <= "000001001011";
rom_data(556) <= "000001001011";
rom_data(557) <= "000001001011";
rom_data(558) <= "000001001100";
rom_data(559) <= "000001001100";
rom_data(560) <= "000001001100";
rom_data(561) <= "000001001100";
rom_data(562) <= "000001001101";
rom_data(563) <= "000001001101";
rom_data(564) <= "000001001101";
rom_data(565) <= "000001001101";
rom_data(566) <= "000001001110";
rom_data(567) <= "000001001110";
rom_data(568) <= "000001001110";
rom_data(569) <= "000001001111";
rom_data(570) <= "000001001111";
rom_data(571) <= "000001001111";
rom_data(572) <= "000001001111";
rom_data(573) <= "000001010000";
rom_data(574) <= "000001010000";
rom_data(575) <= "000001010000";
rom_data(576) <= "000001010001";
rom_data(577) <= "000001010001";
rom_data(578) <= "000001010001";
rom_data(579) <= "000001010001";
rom_data(580) <= "000001010010";
rom_data(581) <= "000001010010";
rom_data(582) <= "000001010010";
rom_data(583) <= "000001010011";
rom_data(584) <= "000001010011";
rom_data(585) <= "000001010011";
rom_data(586) <= "000001010011";
rom_data(587) <= "000001010100";
rom_data(588) <= "000001010100";
rom_data(589) <= "000001010100";
rom_data(590) <= "000001010101";
rom_data(591) <= "000001010101";
rom_data(592) <= "000001010101";
rom_data(593) <= "000001010101";
rom_data(594) <= "000001010110";
rom_data(595) <= "000001010110";
rom_data(596) <= "000001010110";
rom_data(597) <= "000001010111";
rom_data(598) <= "000001010111";
rom_data(599) <= "000001010111";
rom_data(600) <= "000001010111";
rom_data(601) <= "000001011000";
rom_data(602) <= "000001011000";
rom_data(603) <= "000001011000";
rom_data(604) <= "000001011001";
rom_data(605) <= "000001011001";
rom_data(606) <= "000001011001";
rom_data(607) <= "000001011001";
rom_data(608) <= "000001011010";
rom_data(609) <= "000001011010";
rom_data(610) <= "000001011010";
rom_data(611) <= "000001011011";
rom_data(612) <= "000001011011";
rom_data(613) <= "000001011011";
rom_data(614) <= "000001011100";
rom_data(615) <= "000001011100";
rom_data(616) <= "000001011100";
rom_data(617) <= "000001011100";
rom_data(618) <= "000001011101";
rom_data(619) <= "000001011101";
rom_data(620) <= "000001011101";
rom_data(621) <= "000001011110";
rom_data(622) <= "000001011110";
rom_data(623) <= "000001011110";
rom_data(624) <= "000001011111";
rom_data(625) <= "000001011111";
rom_data(626) <= "000001011111";
rom_data(627) <= "000001100000";
rom_data(628) <= "000001100000";
rom_data(629) <= "000001100000";
rom_data(630) <= "000001100000";
rom_data(631) <= "000001100001";
rom_data(632) <= "000001100001";
rom_data(633) <= "000001100001";
rom_data(634) <= "000001100010";
rom_data(635) <= "000001100010";
rom_data(636) <= "000001100010";
rom_data(637) <= "000001100011";
rom_data(638) <= "000001100011";
rom_data(639) <= "000001100011";
rom_data(640) <= "000001100100";
rom_data(641) <= "000001100100";
rom_data(642) <= "000001100100";
rom_data(643) <= "000001100100";
rom_data(644) <= "000001100101";
rom_data(645) <= "000001100101";
rom_data(646) <= "000001100101";
rom_data(647) <= "000001100110";
rom_data(648) <= "000001100110";
rom_data(649) <= "000001100110";
rom_data(650) <= "000001100111";
rom_data(651) <= "000001100111";
rom_data(652) <= "000001100111";
rom_data(653) <= "000001101000";
rom_data(654) <= "000001101000";
rom_data(655) <= "000001101000";
rom_data(656) <= "000001101001";
rom_data(657) <= "000001101001";
rom_data(658) <= "000001101001";
rom_data(659) <= "000001101010";
rom_data(660) <= "000001101010";
rom_data(661) <= "000001101010";
rom_data(662) <= "000001101011";
rom_data(663) <= "000001101011";
rom_data(664) <= "000001101011";
rom_data(665) <= "000001101011";
rom_data(666) <= "000001101100";
rom_data(667) <= "000001101100";
rom_data(668) <= "000001101100";
rom_data(669) <= "000001101101";
rom_data(670) <= "000001101101";
rom_data(671) <= "000001101101";
rom_data(672) <= "000001101110";
rom_data(673) <= "000001101110";
rom_data(674) <= "000001101110";
rom_data(675) <= "000001101111";
rom_data(676) <= "000001101111";
rom_data(677) <= "000001101111";
rom_data(678) <= "000001110000";
rom_data(679) <= "000001110000";
rom_data(680) <= "000001110000";
rom_data(681) <= "000001110001";
rom_data(682) <= "000001110001";
rom_data(683) <= "000001110001";
rom_data(684) <= "000001110010";
rom_data(685) <= "000001110010";
rom_data(686) <= "000001110010";
rom_data(687) <= "000001110011";
rom_data(688) <= "000001110011";
rom_data(689) <= "000001110011";
rom_data(690) <= "000001110100";
rom_data(691) <= "000001110100";
rom_data(692) <= "000001110100";
rom_data(693) <= "000001110101";
rom_data(694) <= "000001110101";
rom_data(695) <= "000001110101";
rom_data(696) <= "000001110110";
rom_data(697) <= "000001110110";
rom_data(698) <= "000001110110";
rom_data(699) <= "000001110111";
rom_data(700) <= "000001110111";
rom_data(701) <= "000001111000";
rom_data(702) <= "000001111000";
rom_data(703) <= "000001111000";
rom_data(704) <= "000001111001";
rom_data(705) <= "000001111001";
rom_data(706) <= "000001111001";
rom_data(707) <= "000001111010";
rom_data(708) <= "000001111010";
rom_data(709) <= "000001111010";
rom_data(710) <= "000001111011";
rom_data(711) <= "000001111011";
rom_data(712) <= "000001111011";
rom_data(713) <= "000001111100";
rom_data(714) <= "000001111100";
rom_data(715) <= "000001111100";
rom_data(716) <= "000001111101";
rom_data(717) <= "000001111101";
rom_data(718) <= "000001111101";
rom_data(719) <= "000001111110";
rom_data(720) <= "000001111110";
rom_data(721) <= "000001111110";
rom_data(722) <= "000001111111";
rom_data(723) <= "000001111111";
rom_data(724) <= "000010000000";
rom_data(725) <= "000010000000";
rom_data(726) <= "000010000000";
rom_data(727) <= "000010000001";
rom_data(728) <= "000010000001";
rom_data(729) <= "000010000001";
rom_data(730) <= "000010000010";
rom_data(731) <= "000010000010";
rom_data(732) <= "000010000010";
rom_data(733) <= "000010000011";
rom_data(734) <= "000010000011";
rom_data(735) <= "000010000011";
rom_data(736) <= "000010000100";
rom_data(737) <= "000010000100";
rom_data(738) <= "000010000101";
rom_data(739) <= "000010000101";
rom_data(740) <= "000010000101";
rom_data(741) <= "000010000110";
rom_data(742) <= "000010000110";
rom_data(743) <= "000010000110";
rom_data(744) <= "000010000111";
rom_data(745) <= "000010000111";
rom_data(746) <= "000010000111";
rom_data(747) <= "000010001000";
rom_data(748) <= "000010001000";
rom_data(749) <= "000010001000";
rom_data(750) <= "000010001001";
rom_data(751) <= "000010001001";
rom_data(752) <= "000010001010";
rom_data(753) <= "000010001010";
rom_data(754) <= "000010001010";
rom_data(755) <= "000010001011";
rom_data(756) <= "000010001011";
rom_data(757) <= "000010001011";
rom_data(758) <= "000010001100";
rom_data(759) <= "000010001100";
rom_data(760) <= "000010001101";
rom_data(761) <= "000010001101";
rom_data(762) <= "000010001101";
rom_data(763) <= "000010001110";
rom_data(764) <= "000010001110";
rom_data(765) <= "000010001110";
rom_data(766) <= "000010001111";
rom_data(767) <= "000010001111";
rom_data(768) <= "000010010000";
rom_data(769) <= "000010010000";
rom_data(770) <= "000010010000";
rom_data(771) <= "000010010001";
rom_data(772) <= "000010010001";
rom_data(773) <= "000010010001";
rom_data(774) <= "000010010010";
rom_data(775) <= "000010010010";
rom_data(776) <= "000010010011";
rom_data(777) <= "000010010011";
rom_data(778) <= "000010010011";
rom_data(779) <= "000010010100";
rom_data(780) <= "000010010100";
rom_data(781) <= "000010010100";
rom_data(782) <= "000010010101";
rom_data(783) <= "000010010101";
rom_data(784) <= "000010010110";
rom_data(785) <= "000010010110";
rom_data(786) <= "000010010110";
rom_data(787) <= "000010010111";
rom_data(788) <= "000010010111";
rom_data(789) <= "000010011000";
rom_data(790) <= "000010011000";
rom_data(791) <= "000010011000";
rom_data(792) <= "000010011001";
rom_data(793) <= "000010011001";
rom_data(794) <= "000010011001";
rom_data(795) <= "000010011010";
rom_data(796) <= "000010011010";
rom_data(797) <= "000010011011";
rom_data(798) <= "000010011011";
rom_data(799) <= "000010011011";
rom_data(800) <= "000010011100";
rom_data(801) <= "000010011100";
rom_data(802) <= "000010011101";
rom_data(803) <= "000010011101";
rom_data(804) <= "000010011101";
rom_data(805) <= "000010011110";
rom_data(806) <= "000010011110";
rom_data(807) <= "000010011111";
rom_data(808) <= "000010011111";
rom_data(809) <= "000010011111";
rom_data(810) <= "000010100000";
rom_data(811) <= "000010100000";
rom_data(812) <= "000010100001";
rom_data(813) <= "000010100001";
rom_data(814) <= "000010100001";
rom_data(815) <= "000010100010";
rom_data(816) <= "000010100010";
rom_data(817) <= "000010100011";
rom_data(818) <= "000010100011";
rom_data(819) <= "000010100011";
rom_data(820) <= "000010100100";
rom_data(821) <= "000010100100";
rom_data(822) <= "000010100101";
rom_data(823) <= "000010100101";
rom_data(824) <= "000010100101";
rom_data(825) <= "000010100110";
rom_data(826) <= "000010100110";
rom_data(827) <= "000010100111";
rom_data(828) <= "000010100111";
rom_data(829) <= "000010100111";
rom_data(830) <= "000010101000";
rom_data(831) <= "000010101000";
rom_data(832) <= "000010101001";
rom_data(833) <= "000010101001";
rom_data(834) <= "000010101001";
rom_data(835) <= "000010101010";
rom_data(836) <= "000010101010";
rom_data(837) <= "000010101011";
rom_data(838) <= "000010101011";
rom_data(839) <= "000010101011";
rom_data(840) <= "000010101100";
rom_data(841) <= "000010101100";
rom_data(842) <= "000010101101";
rom_data(843) <= "000010101101";
rom_data(844) <= "000010101101";
rom_data(845) <= "000010101110";
rom_data(846) <= "000010101110";
rom_data(847) <= "000010101111";
rom_data(848) <= "000010101111";
rom_data(849) <= "000010110000";
rom_data(850) <= "000010110000";
rom_data(851) <= "000010110000";
rom_data(852) <= "000010110001";
rom_data(853) <= "000010110001";
rom_data(854) <= "000010110010";
rom_data(855) <= "000010110010";
rom_data(856) <= "000010110010";
rom_data(857) <= "000010110011";
rom_data(858) <= "000010110011";
rom_data(859) <= "000010110100";
rom_data(860) <= "000010110100";
rom_data(861) <= "000010110101";
rom_data(862) <= "000010110101";
rom_data(863) <= "000010110101";
rom_data(864) <= "000010110110";
rom_data(865) <= "000010110110";
rom_data(866) <= "000010110111";
rom_data(867) <= "000010110111";
rom_data(868) <= "000010110111";
rom_data(869) <= "000010111000";
rom_data(870) <= "000010111000";
rom_data(871) <= "000010111001";
rom_data(872) <= "000010111001";
rom_data(873) <= "000010111010";
rom_data(874) <= "000010111010";
rom_data(875) <= "000010111010";
rom_data(876) <= "000010111011";
rom_data(877) <= "000010111011";
rom_data(878) <= "000010111100";
rom_data(879) <= "000010111100";
rom_data(880) <= "000010111101";
rom_data(881) <= "000010111101";
rom_data(882) <= "000010111101";
rom_data(883) <= "000010111110";
rom_data(884) <= "000010111110";
rom_data(885) <= "000010111111";
rom_data(886) <= "000010111111";
rom_data(887) <= "000011000000";
rom_data(888) <= "000011000000";
rom_data(889) <= "000011000000";
rom_data(890) <= "000011000001";
rom_data(891) <= "000011000001";
rom_data(892) <= "000011000010";
rom_data(893) <= "000011000010";
rom_data(894) <= "000011000011";
rom_data(895) <= "000011000011";
rom_data(896) <= "000011000100";
rom_data(897) <= "000011000100";
rom_data(898) <= "000011000100";
rom_data(899) <= "000011000101";
rom_data(900) <= "000011000101";
rom_data(901) <= "000011000110";
rom_data(902) <= "000011000110";
rom_data(903) <= "000011000111";
rom_data(904) <= "000011000111";
rom_data(905) <= "000011001000";
rom_data(906) <= "000011001000";
rom_data(907) <= "000011001000";
rom_data(908) <= "000011001001";
rom_data(909) <= "000011001001";
rom_data(910) <= "000011001010";
rom_data(911) <= "000011001010";
rom_data(912) <= "000011001011";
rom_data(913) <= "000011001011";
rom_data(914) <= "000011001100";
rom_data(915) <= "000011001100";
rom_data(916) <= "000011001100";
rom_data(917) <= "000011001101";
rom_data(918) <= "000011001101";
rom_data(919) <= "000011001110";
rom_data(920) <= "000011001110";
rom_data(921) <= "000011001111";
rom_data(922) <= "000011001111";
rom_data(923) <= "000011010000";
rom_data(924) <= "000011010000";
rom_data(925) <= "000011010000";
rom_data(926) <= "000011010001";
rom_data(927) <= "000011010001";
rom_data(928) <= "000011010010";
rom_data(929) <= "000011010010";
rom_data(930) <= "000011010011";
rom_data(931) <= "000011010011";
rom_data(932) <= "000011010100";
rom_data(933) <= "000011010100";
rom_data(934) <= "000011010101";
rom_data(935) <= "000011010101";
rom_data(936) <= "000011010101";
rom_data(937) <= "000011010110";
rom_data(938) <= "000011010110";
rom_data(939) <= "000011010111";
rom_data(940) <= "000011010111";
rom_data(941) <= "000011011000";
rom_data(942) <= "000011011000";
rom_data(943) <= "000011011001";
rom_data(944) <= "000011011001";
rom_data(945) <= "000011011010";
rom_data(946) <= "000011011010";
rom_data(947) <= "000011011011";
rom_data(948) <= "000011011011";
rom_data(949) <= "000011011011";
rom_data(950) <= "000011011100";
rom_data(951) <= "000011011100";
rom_data(952) <= "000011011101";
rom_data(953) <= "000011011101";
rom_data(954) <= "000011011110";
rom_data(955) <= "000011011110";
rom_data(956) <= "000011011111";
rom_data(957) <= "000011011111";
rom_data(958) <= "000011100000";
rom_data(959) <= "000011100000";
rom_data(960) <= "000011100001";
rom_data(961) <= "000011100001";
rom_data(962) <= "000011100001";
rom_data(963) <= "000011100010";
rom_data(964) <= "000011100010";
rom_data(965) <= "000011100011";
rom_data(966) <= "000011100011";
rom_data(967) <= "000011100100";
rom_data(968) <= "000011100100";
rom_data(969) <= "000011100101";
rom_data(970) <= "000011100101";
rom_data(971) <= "000011100110";
rom_data(972) <= "000011100110";
rom_data(973) <= "000011100111";
rom_data(974) <= "000011100111";
rom_data(975) <= "000011101000";
rom_data(976) <= "000011101000";
rom_data(977) <= "000011101001";
rom_data(978) <= "000011101001";
rom_data(979) <= "000011101010";
rom_data(980) <= "000011101010";
rom_data(981) <= "000011101011";
rom_data(982) <= "000011101011";
rom_data(983) <= "000011101011";
rom_data(984) <= "000011101100";
rom_data(985) <= "000011101100";
rom_data(986) <= "000011101101";
rom_data(987) <= "000011101101";
rom_data(988) <= "000011101110";
rom_data(989) <= "000011101110";
rom_data(990) <= "000011101111";
rom_data(991) <= "000011101111";
rom_data(992) <= "000011110000";
rom_data(993) <= "000011110000";
rom_data(994) <= "000011110001";
rom_data(995) <= "000011110001";
rom_data(996) <= "000011110010";
rom_data(997) <= "000011110010";
rom_data(998) <= "000011110011";
rom_data(999) <= "000011110011";
rom_data(1000) <= "000011110100";
rom_data(1001) <= "000011110100";
rom_data(1002) <= "000011110101";
rom_data(1003) <= "000011110101";
rom_data(1004) <= "000011110110";
rom_data(1005) <= "000011110110";
rom_data(1006) <= "000011110111";
rom_data(1007) <= "000011110111";
rom_data(1008) <= "000011111000";
rom_data(1009) <= "000011111000";
rom_data(1010) <= "000011111001";
rom_data(1011) <= "000011111001";
rom_data(1012) <= "000011111010";
rom_data(1013) <= "000011111010";
rom_data(1014) <= "000011111011";
rom_data(1015) <= "000011111011";
rom_data(1016) <= "000011111100";
rom_data(1017) <= "000011111100";
rom_data(1018) <= "000011111101";
rom_data(1019) <= "000011111101";
rom_data(1020) <= "000011111110";
rom_data(1021) <= "000011111110";
rom_data(1022) <= "000011111111";
rom_data(1023) <= "000011111111";
rom_data(1024) <= "000100000000";
rom_data(1025) <= "000100000000";
rom_data(1026) <= "000100000001";
rom_data(1027) <= "000100000001";
rom_data(1028) <= "000100000010";
rom_data(1029) <= "000100000010";
rom_data(1030) <= "000100000011";
rom_data(1031) <= "000100000011";
rom_data(1032) <= "000100000100";
rom_data(1033) <= "000100000100";
rom_data(1034) <= "000100000101";
rom_data(1035) <= "000100000101";
rom_data(1036) <= "000100000110";
rom_data(1037) <= "000100000110";
rom_data(1038) <= "000100000111";
rom_data(1039) <= "000100000111";
rom_data(1040) <= "000100001000";
rom_data(1041) <= "000100001000";
rom_data(1042) <= "000100001001";
rom_data(1043) <= "000100001001";
rom_data(1044) <= "000100001010";
rom_data(1045) <= "000100001010";
rom_data(1046) <= "000100001011";
rom_data(1047) <= "000100001011";
rom_data(1048) <= "000100001100";
rom_data(1049) <= "000100001100";
rom_data(1050) <= "000100001101";
rom_data(1051) <= "000100001101";
rom_data(1052) <= "000100001110";
rom_data(1053) <= "000100001110";
rom_data(1054) <= "000100001111";
rom_data(1055) <= "000100001111";
rom_data(1056) <= "000100010000";
rom_data(1057) <= "000100010000";
rom_data(1058) <= "000100010001";
rom_data(1059) <= "000100010001";
rom_data(1060) <= "000100010010";
rom_data(1061) <= "000100010010";
rom_data(1062) <= "000100010011";
rom_data(1063) <= "000100010011";
rom_data(1064) <= "000100010100";
rom_data(1065) <= "000100010100";
rom_data(1066) <= "000100010101";
rom_data(1067) <= "000100010110";
rom_data(1068) <= "000100010110";
rom_data(1069) <= "000100010111";
rom_data(1070) <= "000100010111";
rom_data(1071) <= "000100011000";
rom_data(1072) <= "000100011000";
rom_data(1073) <= "000100011001";
rom_data(1074) <= "000100011001";
rom_data(1075) <= "000100011010";
rom_data(1076) <= "000100011010";
rom_data(1077) <= "000100011011";
rom_data(1078) <= "000100011011";
rom_data(1079) <= "000100011100";
rom_data(1080) <= "000100011100";
rom_data(1081) <= "000100011101";
rom_data(1082) <= "000100011101";
rom_data(1083) <= "000100011110";
rom_data(1084) <= "000100011110";
rom_data(1085) <= "000100011111";
rom_data(1086) <= "000100100000";
rom_data(1087) <= "000100100000";
rom_data(1088) <= "000100100001";
rom_data(1089) <= "000100100001";
rom_data(1090) <= "000100100010";
rom_data(1091) <= "000100100010";
rom_data(1092) <= "000100100011";
rom_data(1093) <= "000100100011";
rom_data(1094) <= "000100100100";
rom_data(1095) <= "000100100100";
rom_data(1096) <= "000100100101";
rom_data(1097) <= "000100100101";
rom_data(1098) <= "000100100110";
rom_data(1099) <= "000100100110";
rom_data(1100) <= "000100100111";
rom_data(1101) <= "000100101000";
rom_data(1102) <= "000100101000";
rom_data(1103) <= "000100101001";
rom_data(1104) <= "000100101001";
rom_data(1105) <= "000100101010";
rom_data(1106) <= "000100101010";
rom_data(1107) <= "000100101011";
rom_data(1108) <= "000100101011";
rom_data(1109) <= "000100101100";
rom_data(1110) <= "000100101100";
rom_data(1111) <= "000100101101";
rom_data(1112) <= "000100101101";
rom_data(1113) <= "000100101110";
rom_data(1114) <= "000100101111";
rom_data(1115) <= "000100101111";
rom_data(1116) <= "000100110000";
rom_data(1117) <= "000100110000";
rom_data(1118) <= "000100110001";
rom_data(1119) <= "000100110001";
rom_data(1120) <= "000100110010";
rom_data(1121) <= "000100110010";
rom_data(1122) <= "000100110011";
rom_data(1123) <= "000100110011";
rom_data(1124) <= "000100110100";
rom_data(1125) <= "000100110101";
rom_data(1126) <= "000100110101";
rom_data(1127) <= "000100110110";
rom_data(1128) <= "000100110110";
rom_data(1129) <= "000100110111";
rom_data(1130) <= "000100110111";
rom_data(1131) <= "000100111000";
rom_data(1132) <= "000100111000";
rom_data(1133) <= "000100111001";
rom_data(1134) <= "000100111010";
rom_data(1135) <= "000100111010";
rom_data(1136) <= "000100111011";
rom_data(1137) <= "000100111011";
rom_data(1138) <= "000100111100";
rom_data(1139) <= "000100111100";
rom_data(1140) <= "000100111101";
rom_data(1141) <= "000100111101";
rom_data(1142) <= "000100111110";
rom_data(1143) <= "000100111111";
rom_data(1144) <= "000100111111";
rom_data(1145) <= "000101000000";
rom_data(1146) <= "000101000000";
rom_data(1147) <= "000101000001";
rom_data(1148) <= "000101000001";
rom_data(1149) <= "000101000010";
rom_data(1150) <= "000101000010";
rom_data(1151) <= "000101000011";
rom_data(1152) <= "000101000100";
rom_data(1153) <= "000101000100";
rom_data(1154) <= "000101000101";
rom_data(1155) <= "000101000101";
rom_data(1156) <= "000101000110";
rom_data(1157) <= "000101000110";
rom_data(1158) <= "000101000111";
rom_data(1159) <= "000101001000";
rom_data(1160) <= "000101001000";
rom_data(1161) <= "000101001001";
rom_data(1162) <= "000101001001";
rom_data(1163) <= "000101001010";
rom_data(1164) <= "000101001010";
rom_data(1165) <= "000101001011";
rom_data(1166) <= "000101001100";
rom_data(1167) <= "000101001100";
rom_data(1168) <= "000101001101";
rom_data(1169) <= "000101001101";
rom_data(1170) <= "000101001110";
rom_data(1171) <= "000101001110";
rom_data(1172) <= "000101001111";
rom_data(1173) <= "000101010000";
rom_data(1174) <= "000101010000";
rom_data(1175) <= "000101010001";
rom_data(1176) <= "000101010001";
rom_data(1177) <= "000101010010";
rom_data(1178) <= "000101010010";
rom_data(1179) <= "000101010011";
rom_data(1180) <= "000101010100";
rom_data(1181) <= "000101010100";
rom_data(1182) <= "000101010101";
rom_data(1183) <= "000101010101";
rom_data(1184) <= "000101010110";
rom_data(1185) <= "000101010110";
rom_data(1186) <= "000101010111";
rom_data(1187) <= "000101011000";
rom_data(1188) <= "000101011000";
rom_data(1189) <= "000101011001";
rom_data(1190) <= "000101011001";
rom_data(1191) <= "000101011010";
rom_data(1192) <= "000101011010";
rom_data(1193) <= "000101011011";
rom_data(1194) <= "000101011100";
rom_data(1195) <= "000101011100";
rom_data(1196) <= "000101011101";
rom_data(1197) <= "000101011101";
rom_data(1198) <= "000101011110";
rom_data(1199) <= "000101011111";
rom_data(1200) <= "000101011111";
rom_data(1201) <= "000101100000";
rom_data(1202) <= "000101100000";
rom_data(1203) <= "000101100001";
rom_data(1204) <= "000101100001";
rom_data(1205) <= "000101100010";
rom_data(1206) <= "000101100011";
rom_data(1207) <= "000101100011";
rom_data(1208) <= "000101100100";
rom_data(1209) <= "000101100100";
rom_data(1210) <= "000101100101";
rom_data(1211) <= "000101100110";
rom_data(1212) <= "000101100110";
rom_data(1213) <= "000101100111";
rom_data(1214) <= "000101100111";
rom_data(1215) <= "000101101000";
rom_data(1216) <= "000101101001";
rom_data(1217) <= "000101101001";
rom_data(1218) <= "000101101010";
rom_data(1219) <= "000101101010";
rom_data(1220) <= "000101101011";
rom_data(1221) <= "000101101100";
rom_data(1222) <= "000101101100";
rom_data(1223) <= "000101101101";
rom_data(1224) <= "000101101101";
rom_data(1225) <= "000101101110";
rom_data(1226) <= "000101101111";
rom_data(1227) <= "000101101111";
rom_data(1228) <= "000101110000";
rom_data(1229) <= "000101110000";
rom_data(1230) <= "000101110001";
rom_data(1231) <= "000101110010";
rom_data(1232) <= "000101110010";
rom_data(1233) <= "000101110011";
rom_data(1234) <= "000101110011";
rom_data(1235) <= "000101110100";
rom_data(1236) <= "000101110101";
rom_data(1237) <= "000101110101";
rom_data(1238) <= "000101110110";
rom_data(1239) <= "000101110110";
rom_data(1240) <= "000101110111";
rom_data(1241) <= "000101111000";
rom_data(1242) <= "000101111000";
rom_data(1243) <= "000101111001";
rom_data(1244) <= "000101111001";
rom_data(1245) <= "000101111010";
rom_data(1246) <= "000101111011";
rom_data(1247) <= "000101111011";
rom_data(1248) <= "000101111100";
rom_data(1249) <= "000101111100";
rom_data(1250) <= "000101111101";
rom_data(1251) <= "000101111110";
rom_data(1252) <= "000101111110";
rom_data(1253) <= "000101111111";
rom_data(1254) <= "000110000000";
rom_data(1255) <= "000110000000";
rom_data(1256) <= "000110000001";
rom_data(1257) <= "000110000001";
rom_data(1258) <= "000110000010";
rom_data(1259) <= "000110000011";
rom_data(1260) <= "000110000011";
rom_data(1261) <= "000110000100";
rom_data(1262) <= "000110000100";
rom_data(1263) <= "000110000101";
rom_data(1264) <= "000110000110";
rom_data(1265) <= "000110000110";
rom_data(1266) <= "000110000111";
rom_data(1267) <= "000110001000";
rom_data(1268) <= "000110001000";
rom_data(1269) <= "000110001001";
rom_data(1270) <= "000110001001";
rom_data(1271) <= "000110001010";
rom_data(1272) <= "000110001011";
rom_data(1273) <= "000110001011";
rom_data(1274) <= "000110001100";
rom_data(1275) <= "000110001100";
rom_data(1276) <= "000110001101";
rom_data(1277) <= "000110001110";
rom_data(1278) <= "000110001110";
rom_data(1279) <= "000110001111";
rom_data(1280) <= "000110010000";
rom_data(1281) <= "000110010000";
rom_data(1282) <= "000110010001";
rom_data(1283) <= "000110010001";
rom_data(1284) <= "000110010010";
rom_data(1285) <= "000110010011";
rom_data(1286) <= "000110010011";
rom_data(1287) <= "000110010100";
rom_data(1288) <= "000110010101";
rom_data(1289) <= "000110010101";
rom_data(1290) <= "000110010110";
rom_data(1291) <= "000110010111";
rom_data(1292) <= "000110010111";
rom_data(1293) <= "000110011000";
rom_data(1294) <= "000110011000";
rom_data(1295) <= "000110011001";
rom_data(1296) <= "000110011010";
rom_data(1297) <= "000110011010";
rom_data(1298) <= "000110011011";
rom_data(1299) <= "000110011100";
rom_data(1300) <= "000110011100";
rom_data(1301) <= "000110011101";
rom_data(1302) <= "000110011101";
rom_data(1303) <= "000110011110";
rom_data(1304) <= "000110011111";
rom_data(1305) <= "000110011111";
rom_data(1306) <= "000110100000";
rom_data(1307) <= "000110100001";
rom_data(1308) <= "000110100001";
rom_data(1309) <= "000110100010";
rom_data(1310) <= "000110100011";
rom_data(1311) <= "000110100011";
rom_data(1312) <= "000110100100";
rom_data(1313) <= "000110100100";
rom_data(1314) <= "000110100101";
rom_data(1315) <= "000110100110";
rom_data(1316) <= "000110100110";
rom_data(1317) <= "000110100111";
rom_data(1318) <= "000110101000";
rom_data(1319) <= "000110101000";
rom_data(1320) <= "000110101001";
rom_data(1321) <= "000110101010";
rom_data(1322) <= "000110101010";
rom_data(1323) <= "000110101011";
rom_data(1324) <= "000110101100";
rom_data(1325) <= "000110101100";
rom_data(1326) <= "000110101101";
rom_data(1327) <= "000110101110";
rom_data(1328) <= "000110101110";
rom_data(1329) <= "000110101111";
rom_data(1330) <= "000110101111";
rom_data(1331) <= "000110110000";
rom_data(1332) <= "000110110001";
rom_data(1333) <= "000110110001";
rom_data(1334) <= "000110110010";
rom_data(1335) <= "000110110011";
rom_data(1336) <= "000110110011";
rom_data(1337) <= "000110110100";
rom_data(1338) <= "000110110101";
rom_data(1339) <= "000110110101";
rom_data(1340) <= "000110110110";
rom_data(1341) <= "000110110111";
rom_data(1342) <= "000110110111";
rom_data(1343) <= "000110111000";
rom_data(1344) <= "000110111001";
rom_data(1345) <= "000110111001";
rom_data(1346) <= "000110111010";
rom_data(1347) <= "000110111011";
rom_data(1348) <= "000110111011";
rom_data(1349) <= "000110111100";
rom_data(1350) <= "000110111101";
rom_data(1351) <= "000110111101";
rom_data(1352) <= "000110111110";
rom_data(1353) <= "000110111111";
rom_data(1354) <= "000110111111";
rom_data(1355) <= "000111000000";
rom_data(1356) <= "000111000001";
rom_data(1357) <= "000111000001";
rom_data(1358) <= "000111000010";
rom_data(1359) <= "000111000011";
rom_data(1360) <= "000111000011";
rom_data(1361) <= "000111000100";
rom_data(1362) <= "000111000101";
rom_data(1363) <= "000111000101";
rom_data(1364) <= "000111000110";
rom_data(1365) <= "000111000111";
rom_data(1366) <= "000111000111";
rom_data(1367) <= "000111001000";
rom_data(1368) <= "000111001001";
rom_data(1369) <= "000111001001";
rom_data(1370) <= "000111001010";
rom_data(1371) <= "000111001011";
rom_data(1372) <= "000111001011";
rom_data(1373) <= "000111001100";
rom_data(1374) <= "000111001101";
rom_data(1375) <= "000111001101";
rom_data(1376) <= "000111001110";
rom_data(1377) <= "000111001111";
rom_data(1378) <= "000111001111";
rom_data(1379) <= "000111010000";
rom_data(1380) <= "000111010001";
rom_data(1381) <= "000111010001";
rom_data(1382) <= "000111010010";
rom_data(1383) <= "000111010011";
rom_data(1384) <= "000111010011";
rom_data(1385) <= "000111010100";
rom_data(1386) <= "000111010101";
rom_data(1387) <= "000111010101";
rom_data(1388) <= "000111010110";
rom_data(1389) <= "000111010111";
rom_data(1390) <= "000111010111";
rom_data(1391) <= "000111011000";
rom_data(1392) <= "000111011001";
rom_data(1393) <= "000111011001";
rom_data(1394) <= "000111011010";
rom_data(1395) <= "000111011011";
rom_data(1396) <= "000111011011";
rom_data(1397) <= "000111011100";
rom_data(1398) <= "000111011101";
rom_data(1399) <= "000111011101";
rom_data(1400) <= "000111011110";
rom_data(1401) <= "000111011111";
rom_data(1402) <= "000111100000";
rom_data(1403) <= "000111100000";
rom_data(1404) <= "000111100001";
rom_data(1405) <= "000111100010";
rom_data(1406) <= "000111100010";
rom_data(1407) <= "000111100011";
rom_data(1408) <= "000111100100";
rom_data(1409) <= "000111100100";
rom_data(1410) <= "000111100101";
rom_data(1411) <= "000111100110";
rom_data(1412) <= "000111100110";
rom_data(1413) <= "000111100111";
rom_data(1414) <= "000111101000";
rom_data(1415) <= "000111101000";
rom_data(1416) <= "000111101001";
rom_data(1417) <= "000111101010";
rom_data(1418) <= "000111101011";
rom_data(1419) <= "000111101011";
rom_data(1420) <= "000111101100";
rom_data(1421) <= "000111101101";
rom_data(1422) <= "000111101101";
rom_data(1423) <= "000111101110";
rom_data(1424) <= "000111101111";
rom_data(1425) <= "000111101111";
rom_data(1426) <= "000111110000";
rom_data(1427) <= "000111110001";
rom_data(1428) <= "000111110001";
rom_data(1429) <= "000111110010";
rom_data(1430) <= "000111110011";
rom_data(1431) <= "000111110100";
rom_data(1432) <= "000111110100";
rom_data(1433) <= "000111110101";
rom_data(1434) <= "000111110110";
rom_data(1435) <= "000111110110";
rom_data(1436) <= "000111110111";
rom_data(1437) <= "000111111000";
rom_data(1438) <= "000111111000";
rom_data(1439) <= "000111111001";
rom_data(1440) <= "000111111010";
rom_data(1441) <= "000111111011";
rom_data(1442) <= "000111111011";
rom_data(1443) <= "000111111100";
rom_data(1444) <= "000111111101";
rom_data(1445) <= "000111111101";
rom_data(1446) <= "000111111110";
rom_data(1447) <= "000111111111";
rom_data(1448) <= "001000000000";
rom_data(1449) <= "001000000000";
rom_data(1450) <= "001000000001";
rom_data(1451) <= "001000000010";
rom_data(1452) <= "001000000010";
rom_data(1453) <= "001000000011";
rom_data(1454) <= "001000000100";
rom_data(1455) <= "001000000100";
rom_data(1456) <= "001000000101";
rom_data(1457) <= "001000000110";
rom_data(1458) <= "001000000111";
rom_data(1459) <= "001000000111";
rom_data(1460) <= "001000001000";
rom_data(1461) <= "001000001001";
rom_data(1462) <= "001000001001";
rom_data(1463) <= "001000001010";
rom_data(1464) <= "001000001011";
rom_data(1465) <= "001000001100";
rom_data(1466) <= "001000001100";
rom_data(1467) <= "001000001101";
rom_data(1468) <= "001000001110";
rom_data(1469) <= "001000001110";
rom_data(1470) <= "001000001111";
rom_data(1471) <= "001000010000";
rom_data(1472) <= "001000010001";
rom_data(1473) <= "001000010001";
rom_data(1474) <= "001000010010";
rom_data(1475) <= "001000010011";
rom_data(1476) <= "001000010100";
rom_data(1477) <= "001000010100";
rom_data(1478) <= "001000010101";
rom_data(1479) <= "001000010110";
rom_data(1480) <= "001000010110";
rom_data(1481) <= "001000010111";
rom_data(1482) <= "001000011000";
rom_data(1483) <= "001000011001";
rom_data(1484) <= "001000011001";
rom_data(1485) <= "001000011010";
rom_data(1486) <= "001000011011";
rom_data(1487) <= "001000011011";
rom_data(1488) <= "001000011100";
rom_data(1489) <= "001000011101";
rom_data(1490) <= "001000011110";
rom_data(1491) <= "001000011110";
rom_data(1492) <= "001000011111";
rom_data(1493) <= "001000100000";
rom_data(1494) <= "001000100001";
rom_data(1495) <= "001000100001";
rom_data(1496) <= "001000100010";
rom_data(1497) <= "001000100011";
rom_data(1498) <= "001000100011";
rom_data(1499) <= "001000100100";
rom_data(1500) <= "001000100101";
rom_data(1501) <= "001000100110";
rom_data(1502) <= "001000100110";
rom_data(1503) <= "001000100111";
rom_data(1504) <= "001000101000";
rom_data(1505) <= "001000101001";
rom_data(1506) <= "001000101001";
rom_data(1507) <= "001000101010";
rom_data(1508) <= "001000101011";
rom_data(1509) <= "001000101100";
rom_data(1510) <= "001000101100";
rom_data(1511) <= "001000101101";
rom_data(1512) <= "001000101110";
rom_data(1513) <= "001000101111";
rom_data(1514) <= "001000101111";
rom_data(1515) <= "001000110000";
rom_data(1516) <= "001000110001";
rom_data(1517) <= "001000110001";
rom_data(1518) <= "001000110010";
rom_data(1519) <= "001000110011";
rom_data(1520) <= "001000110100";
rom_data(1521) <= "001000110100";
rom_data(1522) <= "001000110101";
rom_data(1523) <= "001000110110";
rom_data(1524) <= "001000110111";
rom_data(1525) <= "001000110111";
rom_data(1526) <= "001000111000";
rom_data(1527) <= "001000111001";
rom_data(1528) <= "001000111010";
rom_data(1529) <= "001000111010";
rom_data(1530) <= "001000111011";
rom_data(1531) <= "001000111100";
rom_data(1532) <= "001000111101";
rom_data(1533) <= "001000111101";
rom_data(1534) <= "001000111110";
rom_data(1535) <= "001000111111";
rom_data(1536) <= "001001000000";
rom_data(1537) <= "001001000000";
rom_data(1538) <= "001001000001";
rom_data(1539) <= "001001000010";
rom_data(1540) <= "001001000011";
rom_data(1541) <= "001001000011";
rom_data(1542) <= "001001000100";
rom_data(1543) <= "001001000101";
rom_data(1544) <= "001001000110";
rom_data(1545) <= "001001000110";
rom_data(1546) <= "001001000111";
rom_data(1547) <= "001001001000";
rom_data(1548) <= "001001001001";
rom_data(1549) <= "001001001001";
rom_data(1550) <= "001001001010";
rom_data(1551) <= "001001001011";
rom_data(1552) <= "001001001100";
rom_data(1553) <= "001001001100";
rom_data(1554) <= "001001001101";
rom_data(1555) <= "001001001110";
rom_data(1556) <= "001001001111";
rom_data(1557) <= "001001010000";
rom_data(1558) <= "001001010000";
rom_data(1559) <= "001001010001";
rom_data(1560) <= "001001010010";
rom_data(1561) <= "001001010011";
rom_data(1562) <= "001001010011";
rom_data(1563) <= "001001010100";
rom_data(1564) <= "001001010101";
rom_data(1565) <= "001001010110";
rom_data(1566) <= "001001010110";
rom_data(1567) <= "001001010111";
rom_data(1568) <= "001001011000";
rom_data(1569) <= "001001011001";
rom_data(1570) <= "001001011001";
rom_data(1571) <= "001001011010";
rom_data(1572) <= "001001011011";
rom_data(1573) <= "001001011100";
rom_data(1574) <= "001001011101";
rom_data(1575) <= "001001011101";
rom_data(1576) <= "001001011110";
rom_data(1577) <= "001001011111";
rom_data(1578) <= "001001100000";
rom_data(1579) <= "001001100000";
rom_data(1580) <= "001001100001";
rom_data(1581) <= "001001100010";
rom_data(1582) <= "001001100011";
rom_data(1583) <= "001001100011";
rom_data(1584) <= "001001100100";
rom_data(1585) <= "001001100101";
rom_data(1586) <= "001001100110";
rom_data(1587) <= "001001100111";
rom_data(1588) <= "001001100111";
rom_data(1589) <= "001001101000";
rom_data(1590) <= "001001101001";
rom_data(1591) <= "001001101010";
rom_data(1592) <= "001001101010";
rom_data(1593) <= "001001101011";
rom_data(1594) <= "001001101100";
rom_data(1595) <= "001001101101";
rom_data(1596) <= "001001101110";
rom_data(1597) <= "001001101110";
rom_data(1598) <= "001001101111";
rom_data(1599) <= "001001110000";
rom_data(1600) <= "001001110001";
rom_data(1601) <= "001001110001";
rom_data(1602) <= "001001110010";
rom_data(1603) <= "001001110011";
rom_data(1604) <= "001001110100";
rom_data(1605) <= "001001110101";
rom_data(1606) <= "001001110101";
rom_data(1607) <= "001001110110";
rom_data(1608) <= "001001110111";
rom_data(1609) <= "001001111000";
rom_data(1610) <= "001001111000";
rom_data(1611) <= "001001111001";
rom_data(1612) <= "001001111010";
rom_data(1613) <= "001001111011";
rom_data(1614) <= "001001111100";
rom_data(1615) <= "001001111100";
rom_data(1616) <= "001001111101";
rom_data(1617) <= "001001111110";
rom_data(1618) <= "001001111111";
rom_data(1619) <= "001010000000";
rom_data(1620) <= "001010000000";
rom_data(1621) <= "001010000001";
rom_data(1622) <= "001010000010";
rom_data(1623) <= "001010000011";
rom_data(1624) <= "001010000100";
rom_data(1625) <= "001010000100";
rom_data(1626) <= "001010000101";
rom_data(1627) <= "001010000110";
rom_data(1628) <= "001010000111";
rom_data(1629) <= "001010001000";
rom_data(1630) <= "001010001000";
rom_data(1631) <= "001010001001";
rom_data(1632) <= "001010001010";
rom_data(1633) <= "001010001011";
rom_data(1634) <= "001010001100";
rom_data(1635) <= "001010001100";
rom_data(1636) <= "001010001101";
rom_data(1637) <= "001010001110";
rom_data(1638) <= "001010001111";
rom_data(1639) <= "001010010000";
rom_data(1640) <= "001010010000";
rom_data(1641) <= "001010010001";
rom_data(1642) <= "001010010010";
rom_data(1643) <= "001010010011";
rom_data(1644) <= "001010010100";
rom_data(1645) <= "001010010100";
rom_data(1646) <= "001010010101";
rom_data(1647) <= "001010010110";
rom_data(1648) <= "001010010111";
rom_data(1649) <= "001010011000";
rom_data(1650) <= "001010011000";
rom_data(1651) <= "001010011001";
rom_data(1652) <= "001010011010";
rom_data(1653) <= "001010011011";
rom_data(1654) <= "001010011100";
rom_data(1655) <= "001010011100";
rom_data(1656) <= "001010011101";
rom_data(1657) <= "001010011110";
rom_data(1658) <= "001010011111";
rom_data(1659) <= "001010100000";
rom_data(1660) <= "001010100000";
rom_data(1661) <= "001010100001";
rom_data(1662) <= "001010100010";
rom_data(1663) <= "001010100011";
rom_data(1664) <= "001010100100";
rom_data(1665) <= "001010100100";
rom_data(1666) <= "001010100101";
rom_data(1667) <= "001010100110";
rom_data(1668) <= "001010100111";
rom_data(1669) <= "001010101000";
rom_data(1670) <= "001010101001";
rom_data(1671) <= "001010101001";
rom_data(1672) <= "001010101010";
rom_data(1673) <= "001010101011";
rom_data(1674) <= "001010101100";
rom_data(1675) <= "001010101101";
rom_data(1676) <= "001010101101";
rom_data(1677) <= "001010101110";
rom_data(1678) <= "001010101111";
rom_data(1679) <= "001010110000";
rom_data(1680) <= "001010110001";
rom_data(1681) <= "001010110010";
rom_data(1682) <= "001010110010";
rom_data(1683) <= "001010110011";
rom_data(1684) <= "001010110100";
rom_data(1685) <= "001010110101";
rom_data(1686) <= "001010110110";
rom_data(1687) <= "001010110110";
rom_data(1688) <= "001010110111";
rom_data(1689) <= "001010111000";
rom_data(1690) <= "001010111001";
rom_data(1691) <= "001010111010";
rom_data(1692) <= "001010111011";
rom_data(1693) <= "001010111011";
rom_data(1694) <= "001010111100";
rom_data(1695) <= "001010111101";
rom_data(1696) <= "001010111110";
rom_data(1697) <= "001010111111";
rom_data(1698) <= "001011000000";
rom_data(1699) <= "001011000000";
rom_data(1700) <= "001011000001";
rom_data(1701) <= "001011000010";
rom_data(1702) <= "001011000011";
rom_data(1703) <= "001011000100";
rom_data(1704) <= "001011000101";
rom_data(1705) <= "001011000101";
rom_data(1706) <= "001011000110";
rom_data(1707) <= "001011000111";
rom_data(1708) <= "001011001000";
rom_data(1709) <= "001011001001";
rom_data(1710) <= "001011001010";
rom_data(1711) <= "001011001010";
rom_data(1712) <= "001011001011";
rom_data(1713) <= "001011001100";
rom_data(1714) <= "001011001101";
rom_data(1715) <= "001011001110";
rom_data(1716) <= "001011001111";
rom_data(1717) <= "001011001111";
rom_data(1718) <= "001011010000";
rom_data(1719) <= "001011010001";
rom_data(1720) <= "001011010010";
rom_data(1721) <= "001011010011";
rom_data(1722) <= "001011010100";
rom_data(1723) <= "001011010100";
rom_data(1724) <= "001011010101";
rom_data(1725) <= "001011010110";
rom_data(1726) <= "001011010111";
rom_data(1727) <= "001011011000";
rom_data(1728) <= "001011011001";
rom_data(1729) <= "001011011010";
rom_data(1730) <= "001011011010";
rom_data(1731) <= "001011011011";
rom_data(1732) <= "001011011100";
rom_data(1733) <= "001011011101";
rom_data(1734) <= "001011011110";
rom_data(1735) <= "001011011111";
rom_data(1736) <= "001011011111";
rom_data(1737) <= "001011100000";
rom_data(1738) <= "001011100001";
rom_data(1739) <= "001011100010";
rom_data(1740) <= "001011100011";
rom_data(1741) <= "001011100100";
rom_data(1742) <= "001011100101";
rom_data(1743) <= "001011100101";
rom_data(1744) <= "001011100110";
rom_data(1745) <= "001011100111";
rom_data(1746) <= "001011101000";
rom_data(1747) <= "001011101001";
rom_data(1748) <= "001011101010";
rom_data(1749) <= "001011101011";
rom_data(1750) <= "001011101011";
rom_data(1751) <= "001011101100";
rom_data(1752) <= "001011101101";
rom_data(1753) <= "001011101110";
rom_data(1754) <= "001011101111";
rom_data(1755) <= "001011110000";
rom_data(1756) <= "001011110001";
rom_data(1757) <= "001011110001";
rom_data(1758) <= "001011110010";
rom_data(1759) <= "001011110011";
rom_data(1760) <= "001011110100";
rom_data(1761) <= "001011110101";
rom_data(1762) <= "001011110110";
rom_data(1763) <= "001011110111";
rom_data(1764) <= "001011110111";
rom_data(1765) <= "001011111000";
rom_data(1766) <= "001011111001";
rom_data(1767) <= "001011111010";
rom_data(1768) <= "001011111011";
rom_data(1769) <= "001011111100";
rom_data(1770) <= "001011111101";
rom_data(1771) <= "001011111101";
rom_data(1772) <= "001011111110";
rom_data(1773) <= "001011111111";
rom_data(1774) <= "001100000000";
rom_data(1775) <= "001100000001";
rom_data(1776) <= "001100000010";
rom_data(1777) <= "001100000011";
rom_data(1778) <= "001100000011";
rom_data(1779) <= "001100000100";
rom_data(1780) <= "001100000101";
rom_data(1781) <= "001100000110";
rom_data(1782) <= "001100000111";
rom_data(1783) <= "001100001000";
rom_data(1784) <= "001100001001";
rom_data(1785) <= "001100001010";
rom_data(1786) <= "001100001010";
rom_data(1787) <= "001100001011";
rom_data(1788) <= "001100001100";
rom_data(1789) <= "001100001101";
rom_data(1790) <= "001100001110";
rom_data(1791) <= "001100001111";
rom_data(1792) <= "001100010000";
rom_data(1793) <= "001100010001";
rom_data(1794) <= "001100010001";
rom_data(1795) <= "001100010010";
rom_data(1796) <= "001100010011";
rom_data(1797) <= "001100010100";
rom_data(1798) <= "001100010101";
rom_data(1799) <= "001100010110";
rom_data(1800) <= "001100010111";
rom_data(1801) <= "001100011000";
rom_data(1802) <= "001100011000";
rom_data(1803) <= "001100011001";
rom_data(1804) <= "001100011010";
rom_data(1805) <= "001100011011";
rom_data(1806) <= "001100011100";
rom_data(1807) <= "001100011101";
rom_data(1808) <= "001100011110";
rom_data(1809) <= "001100011111";
rom_data(1810) <= "001100100000";
rom_data(1811) <= "001100100000";
rom_data(1812) <= "001100100001";
rom_data(1813) <= "001100100010";
rom_data(1814) <= "001100100011";
rom_data(1815) <= "001100100100";
rom_data(1816) <= "001100100101";
rom_data(1817) <= "001100100110";
rom_data(1818) <= "001100100111";
rom_data(1819) <= "001100101000";
rom_data(1820) <= "001100101000";
rom_data(1821) <= "001100101001";
rom_data(1822) <= "001100101010";
rom_data(1823) <= "001100101011";
rom_data(1824) <= "001100101100";
rom_data(1825) <= "001100101101";
rom_data(1826) <= "001100101110";
rom_data(1827) <= "001100101111";
rom_data(1828) <= "001100110000";
rom_data(1829) <= "001100110000";
rom_data(1830) <= "001100110001";
rom_data(1831) <= "001100110010";
rom_data(1832) <= "001100110011";
rom_data(1833) <= "001100110100";
rom_data(1834) <= "001100110101";
rom_data(1835) <= "001100110110";
rom_data(1836) <= "001100110111";
rom_data(1837) <= "001100111000";
rom_data(1838) <= "001100111000";
rom_data(1839) <= "001100111001";
rom_data(1840) <= "001100111010";
rom_data(1841) <= "001100111011";
rom_data(1842) <= "001100111100";
rom_data(1843) <= "001100111101";
rom_data(1844) <= "001100111110";
rom_data(1845) <= "001100111111";
rom_data(1846) <= "001101000000";
rom_data(1847) <= "001101000001";
rom_data(1848) <= "001101000001";
rom_data(1849) <= "001101000010";
rom_data(1850) <= "001101000011";
rom_data(1851) <= "001101000100";
rom_data(1852) <= "001101000101";
rom_data(1853) <= "001101000110";
rom_data(1854) <= "001101000111";
rom_data(1855) <= "001101001000";
rom_data(1856) <= "001101001001";
rom_data(1857) <= "001101001010";
rom_data(1858) <= "001101001011";
rom_data(1859) <= "001101001011";
rom_data(1860) <= "001101001100";
rom_data(1861) <= "001101001101";
rom_data(1862) <= "001101001110";
rom_data(1863) <= "001101001111";
rom_data(1864) <= "001101010000";
rom_data(1865) <= "001101010001";
rom_data(1866) <= "001101010010";
rom_data(1867) <= "001101010011";
rom_data(1868) <= "001101010100";
rom_data(1869) <= "001101010101";
rom_data(1870) <= "001101010101";
rom_data(1871) <= "001101010110";
rom_data(1872) <= "001101010111";
rom_data(1873) <= "001101011000";
rom_data(1874) <= "001101011001";
rom_data(1875) <= "001101011010";
rom_data(1876) <= "001101011011";
rom_data(1877) <= "001101011100";
rom_data(1878) <= "001101011101";
rom_data(1879) <= "001101011110";
rom_data(1880) <= "001101011111";
rom_data(1881) <= "001101100000";
rom_data(1882) <= "001101100000";
rom_data(1883) <= "001101100001";
rom_data(1884) <= "001101100010";
rom_data(1885) <= "001101100011";
rom_data(1886) <= "001101100100";
rom_data(1887) <= "001101100101";
rom_data(1888) <= "001101100110";
rom_data(1889) <= "001101100111";
rom_data(1890) <= "001101101000";
rom_data(1891) <= "001101101001";
rom_data(1892) <= "001101101010";
rom_data(1893) <= "001101101011";
rom_data(1894) <= "001101101100";
rom_data(1895) <= "001101101100";
rom_data(1896) <= "001101101101";
rom_data(1897) <= "001101101110";
rom_data(1898) <= "001101101111";
rom_data(1899) <= "001101110000";
rom_data(1900) <= "001101110001";
rom_data(1901) <= "001101110010";
rom_data(1902) <= "001101110011";
rom_data(1903) <= "001101110100";
rom_data(1904) <= "001101110101";
rom_data(1905) <= "001101110110";
rom_data(1906) <= "001101110111";
rom_data(1907) <= "001101111000";
rom_data(1908) <= "001101111001";
rom_data(1909) <= "001101111001";
rom_data(1910) <= "001101111010";
rom_data(1911) <= "001101111011";
rom_data(1912) <= "001101111100";
rom_data(1913) <= "001101111101";
rom_data(1914) <= "001101111110";
rom_data(1915) <= "001101111111";
rom_data(1916) <= "001110000000";
rom_data(1917) <= "001110000001";
rom_data(1918) <= "001110000010";
rom_data(1919) <= "001110000011";
rom_data(1920) <= "001110000100";
rom_data(1921) <= "001110000101";
rom_data(1922) <= "001110000110";
rom_data(1923) <= "001110000111";
rom_data(1924) <= "001110000111";
rom_data(1925) <= "001110001000";
rom_data(1926) <= "001110001001";
rom_data(1927) <= "001110001010";
rom_data(1928) <= "001110001011";
rom_data(1929) <= "001110001100";
rom_data(1930) <= "001110001101";
rom_data(1931) <= "001110001110";
rom_data(1932) <= "001110001111";
rom_data(1933) <= "001110010000";
rom_data(1934) <= "001110010001";
rom_data(1935) <= "001110010010";
rom_data(1936) <= "001110010011";
rom_data(1937) <= "001110010100";
rom_data(1938) <= "001110010101";
rom_data(1939) <= "001110010110";
rom_data(1940) <= "001110010111";
rom_data(1941) <= "001110011000";
rom_data(1942) <= "001110011000";
rom_data(1943) <= "001110011001";
rom_data(1944) <= "001110011010";
rom_data(1945) <= "001110011011";
rom_data(1946) <= "001110011100";
rom_data(1947) <= "001110011101";
rom_data(1948) <= "001110011110";
rom_data(1949) <= "001110011111";
rom_data(1950) <= "001110100000";
rom_data(1951) <= "001110100001";
rom_data(1952) <= "001110100010";
rom_data(1953) <= "001110100011";
rom_data(1954) <= "001110100100";
rom_data(1955) <= "001110100101";
rom_data(1956) <= "001110100110";
rom_data(1957) <= "001110100111";
rom_data(1958) <= "001110101000";
rom_data(1959) <= "001110101001";
rom_data(1960) <= "001110101010";
rom_data(1961) <= "001110101011";
rom_data(1962) <= "001110101100";
rom_data(1963) <= "001110101100";
rom_data(1964) <= "001110101101";
rom_data(1965) <= "001110101110";
rom_data(1966) <= "001110101111";
rom_data(1967) <= "001110110000";
rom_data(1968) <= "001110110001";
rom_data(1969) <= "001110110010";
rom_data(1970) <= "001110110011";
rom_data(1971) <= "001110110100";
rom_data(1972) <= "001110110101";
rom_data(1973) <= "001110110110";
rom_data(1974) <= "001110110111";
rom_data(1975) <= "001110111000";
rom_data(1976) <= "001110111001";
rom_data(1977) <= "001110111010";
rom_data(1978) <= "001110111011";
rom_data(1979) <= "001110111100";
rom_data(1980) <= "001110111101";
rom_data(1981) <= "001110111110";
rom_data(1982) <= "001110111111";
rom_data(1983) <= "001111000000";
rom_data(1984) <= "001111000001";
rom_data(1985) <= "001111000010";
rom_data(1986) <= "001111000011";
rom_data(1987) <= "001111000100";
rom_data(1988) <= "001111000101";
rom_data(1989) <= "001111000110";
rom_data(1990) <= "001111000111";
rom_data(1991) <= "001111001000";
rom_data(1992) <= "001111001001";
rom_data(1993) <= "001111001001";
rom_data(1994) <= "001111001010";
rom_data(1995) <= "001111001011";
rom_data(1996) <= "001111001100";
rom_data(1997) <= "001111001101";
rom_data(1998) <= "001111001110";
rom_data(1999) <= "001111001111";
rom_data(2000) <= "001111010000";
rom_data(2001) <= "001111010001";
rom_data(2002) <= "001111010010";
rom_data(2003) <= "001111010011";
rom_data(2004) <= "001111010100";
rom_data(2005) <= "001111010101";
rom_data(2006) <= "001111010110";
rom_data(2007) <= "001111010111";
rom_data(2008) <= "001111011000";
rom_data(2009) <= "001111011001";
rom_data(2010) <= "001111011010";
rom_data(2011) <= "001111011011";
rom_data(2012) <= "001111011100";
rom_data(2013) <= "001111011101";
rom_data(2014) <= "001111011110";
rom_data(2015) <= "001111011111";
rom_data(2016) <= "001111100000";
rom_data(2017) <= "001111100001";
rom_data(2018) <= "001111100010";
rom_data(2019) <= "001111100011";
rom_data(2020) <= "001111100100";
rom_data(2021) <= "001111100101";
rom_data(2022) <= "001111100110";
rom_data(2023) <= "001111100111";
rom_data(2024) <= "001111101000";
rom_data(2025) <= "001111101001";
rom_data(2026) <= "001111101010";
rom_data(2027) <= "001111101011";
rom_data(2028) <= "001111101100";
rom_data(2029) <= "001111101101";
rom_data(2030) <= "001111101110";
rom_data(2031) <= "001111101111";
rom_data(2032) <= "001111110000";
rom_data(2033) <= "001111110001";
rom_data(2034) <= "001111110010";
rom_data(2035) <= "001111110011";
rom_data(2036) <= "001111110100";
rom_data(2037) <= "001111110101";
rom_data(2038) <= "001111110110";
rom_data(2039) <= "001111110111";
rom_data(2040) <= "001111111000";
rom_data(2041) <= "001111111001";
rom_data(2042) <= "001111111010";
rom_data(2043) <= "001111111011";
rom_data(2044) <= "001111111100";
rom_data(2045) <= "001111111101";
rom_data(2046) <= "001111111110";
rom_data(2047) <= "001111111111";
rom_data(2048) <= "010000000000";
rom_data(2049) <= "010000000001";
rom_data(2050) <= "010000000010";
rom_data(2051) <= "010000000011";
rom_data(2052) <= "010000000100";
rom_data(2053) <= "010000000101";
rom_data(2054) <= "010000000110";
rom_data(2055) <= "010000000111";
rom_data(2056) <= "010000001000";
rom_data(2057) <= "010000001001";
rom_data(2058) <= "010000001010";
rom_data(2059) <= "010000001011";
rom_data(2060) <= "010000001100";
rom_data(2061) <= "010000001101";
rom_data(2062) <= "010000001110";
rom_data(2063) <= "010000001111";
rom_data(2064) <= "010000010000";
rom_data(2065) <= "010000010001";
rom_data(2066) <= "010000010010";
rom_data(2067) <= "010000010011";
rom_data(2068) <= "010000010100";
rom_data(2069) <= "010000010101";
rom_data(2070) <= "010000010110";
rom_data(2071) <= "010000010111";
rom_data(2072) <= "010000011000";
rom_data(2073) <= "010000011001";
rom_data(2074) <= "010000011010";
rom_data(2075) <= "010000011011";
rom_data(2076) <= "010000011100";
rom_data(2077) <= "010000011101";
rom_data(2078) <= "010000011110";
rom_data(2079) <= "010000011111";
rom_data(2080) <= "010000100000";
rom_data(2081) <= "010000100001";
rom_data(2082) <= "010000100010";
rom_data(2083) <= "010000100011";
rom_data(2084) <= "010000100100";
rom_data(2085) <= "010000100101";
rom_data(2086) <= "010000100110";
rom_data(2087) <= "010000100111";
rom_data(2088) <= "010000101000";
rom_data(2089) <= "010000101001";
rom_data(2090) <= "010000101010";
rom_data(2091) <= "010000101011";
rom_data(2092) <= "010000101100";
rom_data(2093) <= "010000101101";
rom_data(2094) <= "010000101110";
rom_data(2095) <= "010000101111";
rom_data(2096) <= "010000110000";
rom_data(2097) <= "010000110001";
rom_data(2098) <= "010000110010";
rom_data(2099) <= "010000110011";
rom_data(2100) <= "010000110100";
rom_data(2101) <= "010000110101";
rom_data(2102) <= "010000110110";
rom_data(2103) <= "010000111000";
rom_data(2104) <= "010000111001";
rom_data(2105) <= "010000111010";
rom_data(2106) <= "010000111011";
rom_data(2107) <= "010000111100";
rom_data(2108) <= "010000111101";
rom_data(2109) <= "010000111110";
rom_data(2110) <= "010000111111";
rom_data(2111) <= "010001000000";
rom_data(2112) <= "010001000001";
rom_data(2113) <= "010001000010";
rom_data(2114) <= "010001000011";
rom_data(2115) <= "010001000100";
rom_data(2116) <= "010001000101";
rom_data(2117) <= "010001000110";
rom_data(2118) <= "010001000111";
rom_data(2119) <= "010001001000";
rom_data(2120) <= "010001001001";
rom_data(2121) <= "010001001010";
rom_data(2122) <= "010001001011";
rom_data(2123) <= "010001001100";
rom_data(2124) <= "010001001101";
rom_data(2125) <= "010001001110";
rom_data(2126) <= "010001001111";
rom_data(2127) <= "010001010000";
rom_data(2128) <= "010001010001";
rom_data(2129) <= "010001010010";
rom_data(2130) <= "010001010011";
rom_data(2131) <= "010001010100";
rom_data(2132) <= "010001010101";
rom_data(2133) <= "010001010111";
rom_data(2134) <= "010001011000";
rom_data(2135) <= "010001011001";
rom_data(2136) <= "010001011010";
rom_data(2137) <= "010001011011";
rom_data(2138) <= "010001011100";
rom_data(2139) <= "010001011101";
rom_data(2140) <= "010001011110";
rom_data(2141) <= "010001011111";
rom_data(2142) <= "010001100000";
rom_data(2143) <= "010001100001";
rom_data(2144) <= "010001100010";
rom_data(2145) <= "010001100011";
rom_data(2146) <= "010001100100";
rom_data(2147) <= "010001100101";
rom_data(2148) <= "010001100110";
rom_data(2149) <= "010001100111";
rom_data(2150) <= "010001101000";
rom_data(2151) <= "010001101001";
rom_data(2152) <= "010001101010";
rom_data(2153) <= "010001101011";
rom_data(2154) <= "010001101101";
rom_data(2155) <= "010001101110";
rom_data(2156) <= "010001101111";
rom_data(2157) <= "010001110000";
rom_data(2158) <= "010001110001";
rom_data(2159) <= "010001110010";
rom_data(2160) <= "010001110011";
rom_data(2161) <= "010001110100";
rom_data(2162) <= "010001110101";
rom_data(2163) <= "010001110110";
rom_data(2164) <= "010001110111";
rom_data(2165) <= "010001111000";
rom_data(2166) <= "010001111001";
rom_data(2167) <= "010001111010";
rom_data(2168) <= "010001111011";
rom_data(2169) <= "010001111100";
rom_data(2170) <= "010001111101";
rom_data(2171) <= "010001111110";
rom_data(2172) <= "010010000000";
rom_data(2173) <= "010010000001";
rom_data(2174) <= "010010000010";
rom_data(2175) <= "010010000011";
rom_data(2176) <= "010010000100";
rom_data(2177) <= "010010000101";
rom_data(2178) <= "010010000110";
rom_data(2179) <= "010010000111";
rom_data(2180) <= "010010001000";
rom_data(2181) <= "010010001001";
rom_data(2182) <= "010010001010";
rom_data(2183) <= "010010001011";
rom_data(2184) <= "010010001100";
rom_data(2185) <= "010010001101";
rom_data(2186) <= "010010001110";
rom_data(2187) <= "010010010000";
rom_data(2188) <= "010010010001";
rom_data(2189) <= "010010010010";
rom_data(2190) <= "010010010011";
rom_data(2191) <= "010010010100";
rom_data(2192) <= "010010010101";
rom_data(2193) <= "010010010110";
rom_data(2194) <= "010010010111";
rom_data(2195) <= "010010011000";
rom_data(2196) <= "010010011001";
rom_data(2197) <= "010010011010";
rom_data(2198) <= "010010011011";
rom_data(2199) <= "010010011100";
rom_data(2200) <= "010010011101";
rom_data(2201) <= "010010011111";
rom_data(2202) <= "010010100000";
rom_data(2203) <= "010010100001";
rom_data(2204) <= "010010100010";
rom_data(2205) <= "010010100011";
rom_data(2206) <= "010010100100";
rom_data(2207) <= "010010100101";
rom_data(2208) <= "010010100110";
rom_data(2209) <= "010010100111";
rom_data(2210) <= "010010101000";
rom_data(2211) <= "010010101001";
rom_data(2212) <= "010010101010";
rom_data(2213) <= "010010101011";
rom_data(2214) <= "010010101101";
rom_data(2215) <= "010010101110";
rom_data(2216) <= "010010101111";
rom_data(2217) <= "010010110000";
rom_data(2218) <= "010010110001";
rom_data(2219) <= "010010110010";
rom_data(2220) <= "010010110011";
rom_data(2221) <= "010010110100";
rom_data(2222) <= "010010110101";
rom_data(2223) <= "010010110110";
rom_data(2224) <= "010010110111";
rom_data(2225) <= "010010111000";
rom_data(2226) <= "010010111010";
rom_data(2227) <= "010010111011";
rom_data(2228) <= "010010111100";
rom_data(2229) <= "010010111101";
rom_data(2230) <= "010010111110";
rom_data(2231) <= "010010111111";
rom_data(2232) <= "010011000000";
rom_data(2233) <= "010011000001";
rom_data(2234) <= "010011000010";
rom_data(2235) <= "010011000011";
rom_data(2236) <= "010011000100";
rom_data(2237) <= "010011000110";
rom_data(2238) <= "010011000111";
rom_data(2239) <= "010011001000";
rom_data(2240) <= "010011001001";
rom_data(2241) <= "010011001010";
rom_data(2242) <= "010011001011";
rom_data(2243) <= "010011001100";
rom_data(2244) <= "010011001101";
rom_data(2245) <= "010011001110";
rom_data(2246) <= "010011001111";
rom_data(2247) <= "010011010000";
rom_data(2248) <= "010011010010";
rom_data(2249) <= "010011010011";
rom_data(2250) <= "010011010100";
rom_data(2251) <= "010011010101";
rom_data(2252) <= "010011010110";
rom_data(2253) <= "010011010111";
rom_data(2254) <= "010011011000";
rom_data(2255) <= "010011011001";
rom_data(2256) <= "010011011010";
rom_data(2257) <= "010011011011";
rom_data(2258) <= "010011011101";
rom_data(2259) <= "010011011110";
rom_data(2260) <= "010011011111";
rom_data(2261) <= "010011100000";
rom_data(2262) <= "010011100001";
rom_data(2263) <= "010011100010";
rom_data(2264) <= "010011100011";
rom_data(2265) <= "010011100100";
rom_data(2266) <= "010011100101";
rom_data(2267) <= "010011100111";
rom_data(2268) <= "010011101000";
rom_data(2269) <= "010011101001";
rom_data(2270) <= "010011101010";
rom_data(2271) <= "010011101011";
rom_data(2272) <= "010011101100";
rom_data(2273) <= "010011101101";
rom_data(2274) <= "010011101110";
rom_data(2275) <= "010011101111";
rom_data(2276) <= "010011110001";
rom_data(2277) <= "010011110010";
rom_data(2278) <= "010011110011";
rom_data(2279) <= "010011110100";
rom_data(2280) <= "010011110101";
rom_data(2281) <= "010011110110";
rom_data(2282) <= "010011110111";
rom_data(2283) <= "010011111000";
rom_data(2284) <= "010011111001";
rom_data(2285) <= "010011111011";
rom_data(2286) <= "010011111100";
rom_data(2287) <= "010011111101";
rom_data(2288) <= "010011111110";
rom_data(2289) <= "010011111111";
rom_data(2290) <= "010100000000";
rom_data(2291) <= "010100000001";
rom_data(2292) <= "010100000010";
rom_data(2293) <= "010100000011";
rom_data(2294) <= "010100000101";
rom_data(2295) <= "010100000110";
rom_data(2296) <= "010100000111";
rom_data(2297) <= "010100001000";
rom_data(2298) <= "010100001001";
rom_data(2299) <= "010100001010";
rom_data(2300) <= "010100001011";
rom_data(2301) <= "010100001100";
rom_data(2302) <= "010100001110";
rom_data(2303) <= "010100001111";
rom_data(2304) <= "010100010000";
rom_data(2305) <= "010100010001";
rom_data(2306) <= "010100010010";
rom_data(2307) <= "010100010011";
rom_data(2308) <= "010100010100";
rom_data(2309) <= "010100010101";
rom_data(2310) <= "010100010111";
rom_data(2311) <= "010100011000";
rom_data(2312) <= "010100011001";
rom_data(2313) <= "010100011010";
rom_data(2314) <= "010100011011";
rom_data(2315) <= "010100011100";
rom_data(2316) <= "010100011101";
rom_data(2317) <= "010100011110";
rom_data(2318) <= "010100100000";
rom_data(2319) <= "010100100001";
rom_data(2320) <= "010100100010";
rom_data(2321) <= "010100100011";
rom_data(2322) <= "010100100100";
rom_data(2323) <= "010100100101";
rom_data(2324) <= "010100100110";
rom_data(2325) <= "010100101000";
rom_data(2326) <= "010100101001";
rom_data(2327) <= "010100101010";
rom_data(2328) <= "010100101011";
rom_data(2329) <= "010100101100";
rom_data(2330) <= "010100101101";
rom_data(2331) <= "010100101110";
rom_data(2332) <= "010100110000";
rom_data(2333) <= "010100110001";
rom_data(2334) <= "010100110010";
rom_data(2335) <= "010100110011";
rom_data(2336) <= "010100110100";
rom_data(2337) <= "010100110101";
rom_data(2338) <= "010100110110";
rom_data(2339) <= "010100111000";
rom_data(2340) <= "010100111001";
rom_data(2341) <= "010100111010";
rom_data(2342) <= "010100111011";
rom_data(2343) <= "010100111100";
rom_data(2344) <= "010100111101";
rom_data(2345) <= "010100111110";
rom_data(2346) <= "010101000000";
rom_data(2347) <= "010101000001";
rom_data(2348) <= "010101000010";
rom_data(2349) <= "010101000011";
rom_data(2350) <= "010101000100";
rom_data(2351) <= "010101000101";
rom_data(2352) <= "010101000110";
rom_data(2353) <= "010101001000";
rom_data(2354) <= "010101001001";
rom_data(2355) <= "010101001010";
rom_data(2356) <= "010101001011";
rom_data(2357) <= "010101001100";
rom_data(2358) <= "010101001101";
rom_data(2359) <= "010101001110";
rom_data(2360) <= "010101010000";
rom_data(2361) <= "010101010001";
rom_data(2362) <= "010101010010";
rom_data(2363) <= "010101010011";
rom_data(2364) <= "010101010100";
rom_data(2365) <= "010101010101";
rom_data(2366) <= "010101010111";
rom_data(2367) <= "010101011000";
rom_data(2368) <= "010101011001";
rom_data(2369) <= "010101011010";
rom_data(2370) <= "010101011011";
rom_data(2371) <= "010101011100";
rom_data(2372) <= "010101011101";
rom_data(2373) <= "010101011111";
rom_data(2374) <= "010101100000";
rom_data(2375) <= "010101100001";
rom_data(2376) <= "010101100010";
rom_data(2377) <= "010101100011";
rom_data(2378) <= "010101100100";
rom_data(2379) <= "010101100110";
rom_data(2380) <= "010101100111";
rom_data(2381) <= "010101101000";
rom_data(2382) <= "010101101001";
rom_data(2383) <= "010101101010";
rom_data(2384) <= "010101101011";
rom_data(2385) <= "010101101101";
rom_data(2386) <= "010101101110";
rom_data(2387) <= "010101101111";
rom_data(2388) <= "010101110000";
rom_data(2389) <= "010101110001";
rom_data(2390) <= "010101110010";
rom_data(2391) <= "010101110100";
rom_data(2392) <= "010101110101";
rom_data(2393) <= "010101110110";
rom_data(2394) <= "010101110111";
rom_data(2395) <= "010101111000";
rom_data(2396) <= "010101111001";
rom_data(2397) <= "010101111011";
rom_data(2398) <= "010101111100";
rom_data(2399) <= "010101111101";
rom_data(2400) <= "010101111110";
rom_data(2401) <= "010101111111";
rom_data(2402) <= "010110000000";
rom_data(2403) <= "010110000010";
rom_data(2404) <= "010110000011";
rom_data(2405) <= "010110000100";
rom_data(2406) <= "010110000101";
rom_data(2407) <= "010110000110";
rom_data(2408) <= "010110000111";
rom_data(2409) <= "010110001001";
rom_data(2410) <= "010110001010";
rom_data(2411) <= "010110001011";
rom_data(2412) <= "010110001100";
rom_data(2413) <= "010110001101";
rom_data(2414) <= "010110001111";
rom_data(2415) <= "010110010000";
rom_data(2416) <= "010110010001";
rom_data(2417) <= "010110010010";
rom_data(2418) <= "010110010011";
rom_data(2419) <= "010110010100";
rom_data(2420) <= "010110010110";
rom_data(2421) <= "010110010111";
rom_data(2422) <= "010110011000";
rom_data(2423) <= "010110011001";
rom_data(2424) <= "010110011010";
rom_data(2425) <= "010110011100";
rom_data(2426) <= "010110011101";
rom_data(2427) <= "010110011110";
rom_data(2428) <= "010110011111";
rom_data(2429) <= "010110100000";
rom_data(2430) <= "010110100001";
rom_data(2431) <= "010110100011";
rom_data(2432) <= "010110100100";
rom_data(2433) <= "010110100101";
rom_data(2434) <= "010110100110";
rom_data(2435) <= "010110100111";
rom_data(2436) <= "010110101001";
rom_data(2437) <= "010110101010";
rom_data(2438) <= "010110101011";
rom_data(2439) <= "010110101100";
rom_data(2440) <= "010110101101";
rom_data(2441) <= "010110101111";
rom_data(2442) <= "010110110000";
rom_data(2443) <= "010110110001";
rom_data(2444) <= "010110110010";
rom_data(2445) <= "010110110011";
rom_data(2446) <= "010110110101";
rom_data(2447) <= "010110110110";
rom_data(2448) <= "010110110111";
rom_data(2449) <= "010110111000";
rom_data(2450) <= "010110111001";
rom_data(2451) <= "010110111011";
rom_data(2452) <= "010110111100";
rom_data(2453) <= "010110111101";
rom_data(2454) <= "010110111110";
rom_data(2455) <= "010110111111";
rom_data(2456) <= "010111000001";
rom_data(2457) <= "010111000010";
rom_data(2458) <= "010111000011";
rom_data(2459) <= "010111000100";
rom_data(2460) <= "010111000101";
rom_data(2461) <= "010111000111";
rom_data(2462) <= "010111001000";
rom_data(2463) <= "010111001001";
rom_data(2464) <= "010111001010";
rom_data(2465) <= "010111001011";
rom_data(2466) <= "010111001101";
rom_data(2467) <= "010111001110";
rom_data(2468) <= "010111001111";
rom_data(2469) <= "010111010000";
rom_data(2470) <= "010111010001";
rom_data(2471) <= "010111010011";
rom_data(2472) <= "010111010100";
rom_data(2473) <= "010111010101";
rom_data(2474) <= "010111010110";
rom_data(2475) <= "010111010111";
rom_data(2476) <= "010111011001";
rom_data(2477) <= "010111011010";
rom_data(2478) <= "010111011011";
rom_data(2479) <= "010111011100";
rom_data(2480) <= "010111011101";
rom_data(2481) <= "010111011111";
rom_data(2482) <= "010111100000";
rom_data(2483) <= "010111100001";
rom_data(2484) <= "010111100010";
rom_data(2485) <= "010111100011";
rom_data(2486) <= "010111100101";
rom_data(2487) <= "010111100110";
rom_data(2488) <= "010111100111";
rom_data(2489) <= "010111101000";
rom_data(2490) <= "010111101010";
rom_data(2491) <= "010111101011";
rom_data(2492) <= "010111101100";
rom_data(2493) <= "010111101101";
rom_data(2494) <= "010111101110";
rom_data(2495) <= "010111110000";
rom_data(2496) <= "010111110001";
rom_data(2497) <= "010111110010";
rom_data(2498) <= "010111110011";
rom_data(2499) <= "010111110101";
rom_data(2500) <= "010111110110";
rom_data(2501) <= "010111110111";
rom_data(2502) <= "010111111000";
rom_data(2503) <= "010111111001";
rom_data(2504) <= "010111111011";
rom_data(2505) <= "010111111100";
rom_data(2506) <= "010111111101";
rom_data(2507) <= "010111111110";
rom_data(2508) <= "011000000000";
rom_data(2509) <= "011000000001";
rom_data(2510) <= "011000000010";
rom_data(2511) <= "011000000011";
rom_data(2512) <= "011000000100";
rom_data(2513) <= "011000000110";
rom_data(2514) <= "011000000111";
rom_data(2515) <= "011000001000";
rom_data(2516) <= "011000001001";
rom_data(2517) <= "011000001011";
rom_data(2518) <= "011000001100";
rom_data(2519) <= "011000001101";
rom_data(2520) <= "011000001110";
rom_data(2521) <= "011000010000";
rom_data(2522) <= "011000010001";
rom_data(2523) <= "011000010010";
rom_data(2524) <= "011000010011";
rom_data(2525) <= "011000010100";
rom_data(2526) <= "011000010110";
rom_data(2527) <= "011000010111";
rom_data(2528) <= "011000011000";
rom_data(2529) <= "011000011001";
rom_data(2530) <= "011000011011";
rom_data(2531) <= "011000011100";
rom_data(2532) <= "011000011101";
rom_data(2533) <= "011000011110";
rom_data(2534) <= "011000100000";
rom_data(2535) <= "011000100001";
rom_data(2536) <= "011000100010";
rom_data(2537) <= "011000100011";
rom_data(2538) <= "011000100101";
rom_data(2539) <= "011000100110";
rom_data(2540) <= "011000100111";
rom_data(2541) <= "011000101000";
rom_data(2542) <= "011000101001";
rom_data(2543) <= "011000101011";
rom_data(2544) <= "011000101100";
rom_data(2545) <= "011000101101";
rom_data(2546) <= "011000101110";
rom_data(2547) <= "011000110000";
rom_data(2548) <= "011000110001";
rom_data(2549) <= "011000110010";
rom_data(2550) <= "011000110011";
rom_data(2551) <= "011000110101";
rom_data(2552) <= "011000110110";
rom_data(2553) <= "011000110111";
rom_data(2554) <= "011000111000";
rom_data(2555) <= "011000111010";
rom_data(2556) <= "011000111011";
rom_data(2557) <= "011000111100";
rom_data(2558) <= "011000111101";
rom_data(2559) <= "011000111111";
rom_data(2560) <= "011001000000";
rom_data(2561) <= "011001000001";
rom_data(2562) <= "011001000010";
rom_data(2563) <= "011001000100";
rom_data(2564) <= "011001000101";
rom_data(2565) <= "011001000110";
rom_data(2566) <= "011001000111";
rom_data(2567) <= "011001001001";
rom_data(2568) <= "011001001010";
rom_data(2569) <= "011001001011";
rom_data(2570) <= "011001001100";
rom_data(2571) <= "011001001110";
rom_data(2572) <= "011001001111";
rom_data(2573) <= "011001010000";
rom_data(2574) <= "011001010001";
rom_data(2575) <= "011001010011";
rom_data(2576) <= "011001010100";
rom_data(2577) <= "011001010101";
rom_data(2578) <= "011001010110";
rom_data(2579) <= "011001011000";
rom_data(2580) <= "011001011001";
rom_data(2581) <= "011001011010";
rom_data(2582) <= "011001011100";
rom_data(2583) <= "011001011101";
rom_data(2584) <= "011001011110";
rom_data(2585) <= "011001011111";
rom_data(2586) <= "011001100001";
rom_data(2587) <= "011001100010";
rom_data(2588) <= "011001100011";
rom_data(2589) <= "011001100100";
rom_data(2590) <= "011001100110";
rom_data(2591) <= "011001100111";
rom_data(2592) <= "011001101000";
rom_data(2593) <= "011001101001";
rom_data(2594) <= "011001101011";
rom_data(2595) <= "011001101100";
rom_data(2596) <= "011001101101";
rom_data(2597) <= "011001101110";
rom_data(2598) <= "011001110000";
rom_data(2599) <= "011001110001";
rom_data(2600) <= "011001110010";
rom_data(2601) <= "011001110100";
rom_data(2602) <= "011001110101";
rom_data(2603) <= "011001110110";
rom_data(2604) <= "011001110111";
rom_data(2605) <= "011001111001";
rom_data(2606) <= "011001111010";
rom_data(2607) <= "011001111011";
rom_data(2608) <= "011001111100";
rom_data(2609) <= "011001111110";
rom_data(2610) <= "011001111111";
rom_data(2611) <= "011010000000";
rom_data(2612) <= "011010000010";
rom_data(2613) <= "011010000011";
rom_data(2614) <= "011010000100";
rom_data(2615) <= "011010000101";
rom_data(2616) <= "011010000111";
rom_data(2617) <= "011010001000";
rom_data(2618) <= "011010001001";
rom_data(2619) <= "011010001011";
rom_data(2620) <= "011010001100";
rom_data(2621) <= "011010001101";
rom_data(2622) <= "011010001110";
rom_data(2623) <= "011010010000";
rom_data(2624) <= "011010010001";
rom_data(2625) <= "011010010010";
rom_data(2626) <= "011010010011";
rom_data(2627) <= "011010010101";
rom_data(2628) <= "011010010110";
rom_data(2629) <= "011010010111";
rom_data(2630) <= "011010011001";
rom_data(2631) <= "011010011010";
rom_data(2632) <= "011010011011";
rom_data(2633) <= "011010011100";
rom_data(2634) <= "011010011110";
rom_data(2635) <= "011010011111";
rom_data(2636) <= "011010100000";
rom_data(2637) <= "011010100010";
rom_data(2638) <= "011010100011";
rom_data(2639) <= "011010100100";
rom_data(2640) <= "011010100101";
rom_data(2641) <= "011010100111";
rom_data(2642) <= "011010101000";
rom_data(2643) <= "011010101001";
rom_data(2644) <= "011010101011";
rom_data(2645) <= "011010101100";
rom_data(2646) <= "011010101101";
rom_data(2647) <= "011010101111";
rom_data(2648) <= "011010110000";
rom_data(2649) <= "011010110001";
rom_data(2650) <= "011010110010";
rom_data(2651) <= "011010110100";
rom_data(2652) <= "011010110101";
rom_data(2653) <= "011010110110";
rom_data(2654) <= "011010111000";
rom_data(2655) <= "011010111001";
rom_data(2656) <= "011010111010";
rom_data(2657) <= "011010111011";
rom_data(2658) <= "011010111101";
rom_data(2659) <= "011010111110";
rom_data(2660) <= "011010111111";
rom_data(2661) <= "011011000001";
rom_data(2662) <= "011011000010";
rom_data(2663) <= "011011000011";
rom_data(2664) <= "011011000101";
rom_data(2665) <= "011011000110";
rom_data(2666) <= "011011000111";
rom_data(2667) <= "011011001000";
rom_data(2668) <= "011011001010";
rom_data(2669) <= "011011001011";
rom_data(2670) <= "011011001100";
rom_data(2671) <= "011011001110";
rom_data(2672) <= "011011001111";
rom_data(2673) <= "011011010000";
rom_data(2674) <= "011011010010";
rom_data(2675) <= "011011010011";
rom_data(2676) <= "011011010100";
rom_data(2677) <= "011011010110";
rom_data(2678) <= "011011010111";
rom_data(2679) <= "011011011000";
rom_data(2680) <= "011011011001";
rom_data(2681) <= "011011011011";
rom_data(2682) <= "011011011100";
rom_data(2683) <= "011011011101";
rom_data(2684) <= "011011011111";
rom_data(2685) <= "011011100000";
rom_data(2686) <= "011011100001";
rom_data(2687) <= "011011100011";
rom_data(2688) <= "011011100100";
rom_data(2689) <= "011011100101";
rom_data(2690) <= "011011100111";
rom_data(2691) <= "011011101000";
rom_data(2692) <= "011011101001";
rom_data(2693) <= "011011101011";
rom_data(2694) <= "011011101100";
rom_data(2695) <= "011011101101";
rom_data(2696) <= "011011101110";
rom_data(2697) <= "011011110000";
rom_data(2698) <= "011011110001";
rom_data(2699) <= "011011110010";
rom_data(2700) <= "011011110100";
rom_data(2701) <= "011011110101";
rom_data(2702) <= "011011110110";
rom_data(2703) <= "011011111000";
rom_data(2704) <= "011011111001";
rom_data(2705) <= "011011111010";
rom_data(2706) <= "011011111100";
rom_data(2707) <= "011011111101";
rom_data(2708) <= "011011111110";
rom_data(2709) <= "011100000000";
rom_data(2710) <= "011100000001";
rom_data(2711) <= "011100000010";
rom_data(2712) <= "011100000100";
rom_data(2713) <= "011100000101";
rom_data(2714) <= "011100000110";
rom_data(2715) <= "011100001000";
rom_data(2716) <= "011100001001";
rom_data(2717) <= "011100001010";
rom_data(2718) <= "011100001100";
rom_data(2719) <= "011100001101";
rom_data(2720) <= "011100001110";
rom_data(2721) <= "011100010000";
rom_data(2722) <= "011100010001";
rom_data(2723) <= "011100010010";
rom_data(2724) <= "011100010100";
rom_data(2725) <= "011100010101";
rom_data(2726) <= "011100010110";
rom_data(2727) <= "011100011000";
rom_data(2728) <= "011100011001";
rom_data(2729) <= "011100011010";
rom_data(2730) <= "011100011100";
rom_data(2731) <= "011100011101";
rom_data(2732) <= "011100011110";
rom_data(2733) <= "011100100000";
rom_data(2734) <= "011100100001";
rom_data(2735) <= "011100100010";
rom_data(2736) <= "011100100100";
rom_data(2737) <= "011100100101";
rom_data(2738) <= "011100100110";
rom_data(2739) <= "011100101000";
rom_data(2740) <= "011100101001";
rom_data(2741) <= "011100101010";
rom_data(2742) <= "011100101100";
rom_data(2743) <= "011100101101";
rom_data(2744) <= "011100101110";
rom_data(2745) <= "011100110000";
rom_data(2746) <= "011100110001";
rom_data(2747) <= "011100110010";
rom_data(2748) <= "011100110100";
rom_data(2749) <= "011100110101";
rom_data(2750) <= "011100110110";
rom_data(2751) <= "011100111000";
rom_data(2752) <= "011100111001";
rom_data(2753) <= "011100111010";
rom_data(2754) <= "011100111100";
rom_data(2755) <= "011100111101";
rom_data(2756) <= "011100111110";
rom_data(2757) <= "011101000000";
rom_data(2758) <= "011101000001";
rom_data(2759) <= "011101000010";
rom_data(2760) <= "011101000100";
rom_data(2761) <= "011101000101";
rom_data(2762) <= "011101000110";
rom_data(2763) <= "011101001000";
rom_data(2764) <= "011101001001";
rom_data(2765) <= "011101001010";
rom_data(2766) <= "011101001100";
rom_data(2767) <= "011101001101";
rom_data(2768) <= "011101001111";
rom_data(2769) <= "011101010000";
rom_data(2770) <= "011101010001";
rom_data(2771) <= "011101010011";
rom_data(2772) <= "011101010100";
rom_data(2773) <= "011101010101";
rom_data(2774) <= "011101010111";
rom_data(2775) <= "011101011000";
rom_data(2776) <= "011101011001";
rom_data(2777) <= "011101011011";
rom_data(2778) <= "011101011100";
rom_data(2779) <= "011101011101";
rom_data(2780) <= "011101011111";
rom_data(2781) <= "011101100000";
rom_data(2782) <= "011101100001";
rom_data(2783) <= "011101100011";
rom_data(2784) <= "011101100100";
rom_data(2785) <= "011101100110";
rom_data(2786) <= "011101100111";
rom_data(2787) <= "011101101000";
rom_data(2788) <= "011101101010";
rom_data(2789) <= "011101101011";
rom_data(2790) <= "011101101100";
rom_data(2791) <= "011101101110";
rom_data(2792) <= "011101101111";
rom_data(2793) <= "011101110000";
rom_data(2794) <= "011101110010";
rom_data(2795) <= "011101110011";
rom_data(2796) <= "011101110101";
rom_data(2797) <= "011101110110";
rom_data(2798) <= "011101110111";
rom_data(2799) <= "011101111001";
rom_data(2800) <= "011101111010";
rom_data(2801) <= "011101111011";
rom_data(2802) <= "011101111101";
rom_data(2803) <= "011101111110";
rom_data(2804) <= "011110000000";
rom_data(2805) <= "011110000001";
rom_data(2806) <= "011110000010";
rom_data(2807) <= "011110000100";
rom_data(2808) <= "011110000101";
rom_data(2809) <= "011110000110";
rom_data(2810) <= "011110001000";
rom_data(2811) <= "011110001001";
rom_data(2812) <= "011110001010";
rom_data(2813) <= "011110001100";
rom_data(2814) <= "011110001101";
rom_data(2815) <= "011110001111";
rom_data(2816) <= "011110010000";
rom_data(2817) <= "011110010001";
rom_data(2818) <= "011110010011";
rom_data(2819) <= "011110010100";
rom_data(2820) <= "011110010101";
rom_data(2821) <= "011110010111";
rom_data(2822) <= "011110011000";
rom_data(2823) <= "011110011010";
rom_data(2824) <= "011110011011";
rom_data(2825) <= "011110011100";
rom_data(2826) <= "011110011110";
rom_data(2827) <= "011110011111";
rom_data(2828) <= "011110100001";
rom_data(2829) <= "011110100010";
rom_data(2830) <= "011110100011";
rom_data(2831) <= "011110100101";
rom_data(2832) <= "011110100110";
rom_data(2833) <= "011110100111";
rom_data(2834) <= "011110101001";
rom_data(2835) <= "011110101010";
rom_data(2836) <= "011110101100";
rom_data(2837) <= "011110101101";
rom_data(2838) <= "011110101110";
rom_data(2839) <= "011110110000";
rom_data(2840) <= "011110110001";
rom_data(2841) <= "011110110011";
rom_data(2842) <= "011110110100";
rom_data(2843) <= "011110110101";
rom_data(2844) <= "011110110111";
rom_data(2845) <= "011110111000";
rom_data(2846) <= "011110111001";
rom_data(2847) <= "011110111011";
rom_data(2848) <= "011110111100";
rom_data(2849) <= "011110111110";
rom_data(2850) <= "011110111111";
rom_data(2851) <= "011111000000";
rom_data(2852) <= "011111000010";
rom_data(2853) <= "011111000011";
rom_data(2854) <= "011111000101";
rom_data(2855) <= "011111000110";
rom_data(2856) <= "011111000111";
rom_data(2857) <= "011111001001";
rom_data(2858) <= "011111001010";
rom_data(2859) <= "011111001100";
rom_data(2860) <= "011111001101";
rom_data(2861) <= "011111001110";
rom_data(2862) <= "011111010000";
rom_data(2863) <= "011111010001";
rom_data(2864) <= "011111010011";
rom_data(2865) <= "011111010100";
rom_data(2866) <= "011111010101";
rom_data(2867) <= "011111010111";
rom_data(2868) <= "011111011000";
rom_data(2869) <= "011111011010";
rom_data(2870) <= "011111011011";
rom_data(2871) <= "011111011100";
rom_data(2872) <= "011111011110";
rom_data(2873) <= "011111011111";
rom_data(2874) <= "011111100001";
rom_data(2875) <= "011111100010";
rom_data(2876) <= "011111100011";
rom_data(2877) <= "011111100101";
rom_data(2878) <= "011111100110";
rom_data(2879) <= "011111101000";
rom_data(2880) <= "011111101001";
rom_data(2881) <= "011111101010";
rom_data(2882) <= "011111101100";
rom_data(2883) <= "011111101101";
rom_data(2884) <= "011111101111";
rom_data(2885) <= "011111110000";
rom_data(2886) <= "011111110001";
rom_data(2887) <= "011111110011";
rom_data(2888) <= "011111110100";
rom_data(2889) <= "011111110110";
rom_data(2890) <= "011111110111";
rom_data(2891) <= "011111111000";
rom_data(2892) <= "011111111010";
rom_data(2893) <= "011111111011";
rom_data(2894) <= "011111111101";
rom_data(2895) <= "011111111110";
rom_data(2896) <= "100000000000";
rom_data(2897) <= "100000000001";
rom_data(2898) <= "100000000010";
rom_data(2899) <= "100000000100";
rom_data(2900) <= "100000000101";
rom_data(2901) <= "100000000111";
rom_data(2902) <= "100000001000";
rom_data(2903) <= "100000001001";
rom_data(2904) <= "100000001011";
rom_data(2905) <= "100000001100";
rom_data(2906) <= "100000001110";
rom_data(2907) <= "100000001111";
rom_data(2908) <= "100000010001";
rom_data(2909) <= "100000010010";
rom_data(2910) <= "100000010011";
rom_data(2911) <= "100000010101";
rom_data(2912) <= "100000010110";
rom_data(2913) <= "100000011000";
rom_data(2914) <= "100000011001";
rom_data(2915) <= "100000011011";
rom_data(2916) <= "100000011100";
rom_data(2917) <= "100000011101";
rom_data(2918) <= "100000011111";
rom_data(2919) <= "100000100000";
rom_data(2920) <= "100000100010";
rom_data(2921) <= "100000100011";
rom_data(2922) <= "100000100101";
rom_data(2923) <= "100000100110";
rom_data(2924) <= "100000100111";
rom_data(2925) <= "100000101001";
rom_data(2926) <= "100000101010";
rom_data(2927) <= "100000101100";
rom_data(2928) <= "100000101101";
rom_data(2929) <= "100000101111";
rom_data(2930) <= "100000110000";
rom_data(2931) <= "100000110001";
rom_data(2932) <= "100000110011";
rom_data(2933) <= "100000110100";
rom_data(2934) <= "100000110110";
rom_data(2935) <= "100000110111";
rom_data(2936) <= "100000111001";
rom_data(2937) <= "100000111010";
rom_data(2938) <= "100000111011";
rom_data(2939) <= "100000111101";
rom_data(2940) <= "100000111110";
rom_data(2941) <= "100001000000";
rom_data(2942) <= "100001000001";
rom_data(2943) <= "100001000011";
rom_data(2944) <= "100001000100";
rom_data(2945) <= "100001000101";
rom_data(2946) <= "100001000111";
rom_data(2947) <= "100001001000";
rom_data(2948) <= "100001001010";
rom_data(2949) <= "100001001011";
rom_data(2950) <= "100001001101";
rom_data(2951) <= "100001001110";
rom_data(2952) <= "100001010000";
rom_data(2953) <= "100001010001";
rom_data(2954) <= "100001010010";
rom_data(2955) <= "100001010100";
rom_data(2956) <= "100001010101";
rom_data(2957) <= "100001010111";
rom_data(2958) <= "100001011000";
rom_data(2959) <= "100001011010";
rom_data(2960) <= "100001011011";
rom_data(2961) <= "100001011101";
rom_data(2962) <= "100001011110";
rom_data(2963) <= "100001011111";
rom_data(2964) <= "100001100001";
rom_data(2965) <= "100001100010";
rom_data(2966) <= "100001100100";
rom_data(2967) <= "100001100101";
rom_data(2968) <= "100001100111";
rom_data(2969) <= "100001101000";
rom_data(2970) <= "100001101010";
rom_data(2971) <= "100001101011";
rom_data(2972) <= "100001101100";
rom_data(2973) <= "100001101110";
rom_data(2974) <= "100001101111";
rom_data(2975) <= "100001110001";
rom_data(2976) <= "100001110010";
rom_data(2977) <= "100001110100";
rom_data(2978) <= "100001110101";
rom_data(2979) <= "100001110111";
rom_data(2980) <= "100001111000";
rom_data(2981) <= "100001111010";
rom_data(2982) <= "100001111011";
rom_data(2983) <= "100001111100";
rom_data(2984) <= "100001111110";
rom_data(2985) <= "100001111111";
rom_data(2986) <= "100010000001";
rom_data(2987) <= "100010000010";
rom_data(2988) <= "100010000100";
rom_data(2989) <= "100010000101";
rom_data(2990) <= "100010000111";
rom_data(2991) <= "100010001000";
rom_data(2992) <= "100010001010";
rom_data(2993) <= "100010001011";
rom_data(2994) <= "100010001101";
rom_data(2995) <= "100010001110";
rom_data(2996) <= "100010001111";
rom_data(2997) <= "100010010001";
rom_data(2998) <= "100010010010";
rom_data(2999) <= "100010010100";
rom_data(3000) <= "100010010101";
rom_data(3001) <= "100010010111";
rom_data(3002) <= "100010011000";
rom_data(3003) <= "100010011010";
rom_data(3004) <= "100010011011";
rom_data(3005) <= "100010011101";
rom_data(3006) <= "100010011110";
rom_data(3007) <= "100010100000";
rom_data(3008) <= "100010100001";
rom_data(3009) <= "100010100011";
rom_data(3010) <= "100010100100";
rom_data(3011) <= "100010100101";
rom_data(3012) <= "100010100111";
rom_data(3013) <= "100010101000";
rom_data(3014) <= "100010101010";
rom_data(3015) <= "100010101011";
rom_data(3016) <= "100010101101";
rom_data(3017) <= "100010101110";
rom_data(3018) <= "100010110000";
rom_data(3019) <= "100010110001";
rom_data(3020) <= "100010110011";
rom_data(3021) <= "100010110100";
rom_data(3022) <= "100010110110";
rom_data(3023) <= "100010110111";
rom_data(3024) <= "100010111001";
rom_data(3025) <= "100010111010";
rom_data(3026) <= "100010111100";
rom_data(3027) <= "100010111101";
rom_data(3028) <= "100010111111";
rom_data(3029) <= "100011000000";
rom_data(3030) <= "100011000001";
rom_data(3031) <= "100011000011";
rom_data(3032) <= "100011000100";
rom_data(3033) <= "100011000110";
rom_data(3034) <= "100011000111";
rom_data(3035) <= "100011001001";
rom_data(3036) <= "100011001010";
rom_data(3037) <= "100011001100";
rom_data(3038) <= "100011001101";
rom_data(3039) <= "100011001111";
rom_data(3040) <= "100011010000";
rom_data(3041) <= "100011010010";
rom_data(3042) <= "100011010011";
rom_data(3043) <= "100011010101";
rom_data(3044) <= "100011010110";
rom_data(3045) <= "100011011000";
rom_data(3046) <= "100011011001";
rom_data(3047) <= "100011011011";
rom_data(3048) <= "100011011100";
rom_data(3049) <= "100011011110";
rom_data(3050) <= "100011011111";
rom_data(3051) <= "100011100001";
rom_data(3052) <= "100011100010";
rom_data(3053) <= "100011100100";
rom_data(3054) <= "100011100101";
rom_data(3055) <= "100011100111";
rom_data(3056) <= "100011101000";
rom_data(3057) <= "100011101010";
rom_data(3058) <= "100011101011";
rom_data(3059) <= "100011101101";
rom_data(3060) <= "100011101110";
rom_data(3061) <= "100011110000";
rom_data(3062) <= "100011110001";
rom_data(3063) <= "100011110011";
rom_data(3064) <= "100011110100";
rom_data(3065) <= "100011110110";
rom_data(3066) <= "100011110111";
rom_data(3067) <= "100011111001";
rom_data(3068) <= "100011111010";
rom_data(3069) <= "100011111100";
rom_data(3070) <= "100011111101";
rom_data(3071) <= "100011111111";
rom_data(3072) <= "100100000000";
rom_data(3073) <= "100100000010";
rom_data(3074) <= "100100000011";
rom_data(3075) <= "100100000101";
rom_data(3076) <= "100100000110";
rom_data(3077) <= "100100001000";
rom_data(3078) <= "100100001001";
rom_data(3079) <= "100100001011";
rom_data(3080) <= "100100001100";
rom_data(3081) <= "100100001110";
rom_data(3082) <= "100100001111";
rom_data(3083) <= "100100010001";
rom_data(3084) <= "100100010010";
rom_data(3085) <= "100100010100";
rom_data(3086) <= "100100010101";
rom_data(3087) <= "100100010111";
rom_data(3088) <= "100100011000";
rom_data(3089) <= "100100011010";
rom_data(3090) <= "100100011011";
rom_data(3091) <= "100100011101";
rom_data(3092) <= "100100011110";
rom_data(3093) <= "100100100000";
rom_data(3094) <= "100100100001";
rom_data(3095) <= "100100100011";
rom_data(3096) <= "100100100100";
rom_data(3097) <= "100100100110";
rom_data(3098) <= "100100100111";
rom_data(3099) <= "100100101001";
rom_data(3100) <= "100100101010";
rom_data(3101) <= "100100101100";
rom_data(3102) <= "100100101101";
rom_data(3103) <= "100100101111";
rom_data(3104) <= "100100110000";
rom_data(3105) <= "100100110010";
rom_data(3106) <= "100100110011";
rom_data(3107) <= "100100110101";
rom_data(3108) <= "100100110110";
rom_data(3109) <= "100100111000";
rom_data(3110) <= "100100111001";
rom_data(3111) <= "100100111011";
rom_data(3112) <= "100100111100";
rom_data(3113) <= "100100111110";
rom_data(3114) <= "100101000000";
rom_data(3115) <= "100101000001";
rom_data(3116) <= "100101000011";
rom_data(3117) <= "100101000100";
rom_data(3118) <= "100101000110";
rom_data(3119) <= "100101000111";
rom_data(3120) <= "100101001001";
rom_data(3121) <= "100101001010";
rom_data(3122) <= "100101001100";
rom_data(3123) <= "100101001101";
rom_data(3124) <= "100101001111";
rom_data(3125) <= "100101010000";
rom_data(3126) <= "100101010010";
rom_data(3127) <= "100101010011";
rom_data(3128) <= "100101010101";
rom_data(3129) <= "100101010110";
rom_data(3130) <= "100101011000";
rom_data(3131) <= "100101011001";
rom_data(3132) <= "100101011011";
rom_data(3133) <= "100101011100";
rom_data(3134) <= "100101011110";
rom_data(3135) <= "100101100000";
rom_data(3136) <= "100101100001";
rom_data(3137) <= "100101100011";
rom_data(3138) <= "100101100100";
rom_data(3139) <= "100101100110";
rom_data(3140) <= "100101100111";
rom_data(3141) <= "100101101001";
rom_data(3142) <= "100101101010";
rom_data(3143) <= "100101101100";
rom_data(3144) <= "100101101101";
rom_data(3145) <= "100101101111";
rom_data(3146) <= "100101110000";
rom_data(3147) <= "100101110010";
rom_data(3148) <= "100101110100";
rom_data(3149) <= "100101110101";
rom_data(3150) <= "100101110111";
rom_data(3151) <= "100101111000";
rom_data(3152) <= "100101111010";
rom_data(3153) <= "100101111011";
rom_data(3154) <= "100101111101";
rom_data(3155) <= "100101111110";
rom_data(3156) <= "100110000000";
rom_data(3157) <= "100110000001";
rom_data(3158) <= "100110000011";
rom_data(3159) <= "100110000100";
rom_data(3160) <= "100110000110";
rom_data(3161) <= "100110001000";
rom_data(3162) <= "100110001001";
rom_data(3163) <= "100110001011";
rom_data(3164) <= "100110001100";
rom_data(3165) <= "100110001110";
rom_data(3166) <= "100110001111";
rom_data(3167) <= "100110010001";
rom_data(3168) <= "100110010010";
rom_data(3169) <= "100110010100";
rom_data(3170) <= "100110010101";
rom_data(3171) <= "100110010111";
rom_data(3172) <= "100110011001";
rom_data(3173) <= "100110011010";
rom_data(3174) <= "100110011100";
rom_data(3175) <= "100110011101";
rom_data(3176) <= "100110011111";
rom_data(3177) <= "100110100000";
rom_data(3178) <= "100110100010";
rom_data(3179) <= "100110100011";
rom_data(3180) <= "100110100101";
rom_data(3181) <= "100110100111";
rom_data(3182) <= "100110101000";
rom_data(3183) <= "100110101010";
rom_data(3184) <= "100110101011";
rom_data(3185) <= "100110101101";
rom_data(3186) <= "100110101110";
rom_data(3187) <= "100110110000";
rom_data(3188) <= "100110110001";
rom_data(3189) <= "100110110011";
rom_data(3190) <= "100110110101";
rom_data(3191) <= "100110110110";
rom_data(3192) <= "100110111000";
rom_data(3193) <= "100110111001";
rom_data(3194) <= "100110111011";
rom_data(3195) <= "100110111100";
rom_data(3196) <= "100110111110";
rom_data(3197) <= "100110111111";
rom_data(3198) <= "100111000001";
rom_data(3199) <= "100111000011";
rom_data(3200) <= "100111000100";
rom_data(3201) <= "100111000110";
rom_data(3202) <= "100111000111";
rom_data(3203) <= "100111001001";
rom_data(3204) <= "100111001010";
rom_data(3205) <= "100111001100";
rom_data(3206) <= "100111001101";
rom_data(3207) <= "100111001111";
rom_data(3208) <= "100111010001";
rom_data(3209) <= "100111010010";
rom_data(3210) <= "100111010100";
rom_data(3211) <= "100111010101";
rom_data(3212) <= "100111010111";
rom_data(3213) <= "100111011000";
rom_data(3214) <= "100111011010";
rom_data(3215) <= "100111011100";
rom_data(3216) <= "100111011101";
rom_data(3217) <= "100111011111";
rom_data(3218) <= "100111100000";
rom_data(3219) <= "100111100010";
rom_data(3220) <= "100111100011";
rom_data(3221) <= "100111100101";
rom_data(3222) <= "100111100111";
rom_data(3223) <= "100111101000";
rom_data(3224) <= "100111101010";
rom_data(3225) <= "100111101011";
rom_data(3226) <= "100111101101";
rom_data(3227) <= "100111101110";
rom_data(3228) <= "100111110000";
rom_data(3229) <= "100111110010";
rom_data(3230) <= "100111110011";
rom_data(3231) <= "100111110101";
rom_data(3232) <= "100111110110";
rom_data(3233) <= "100111111000";
rom_data(3234) <= "100111111010";
rom_data(3235) <= "100111111011";
rom_data(3236) <= "100111111101";
rom_data(3237) <= "100111111110";
rom_data(3238) <= "101000000000";
rom_data(3239) <= "101000000001";
rom_data(3240) <= "101000000011";
rom_data(3241) <= "101000000101";
rom_data(3242) <= "101000000110";
rom_data(3243) <= "101000001000";
rom_data(3244) <= "101000001001";
rom_data(3245) <= "101000001011";
rom_data(3246) <= "101000001101";
rom_data(3247) <= "101000001110";
rom_data(3248) <= "101000010000";
rom_data(3249) <= "101000010001";
rom_data(3250) <= "101000010011";
rom_data(3251) <= "101000010100";
rom_data(3252) <= "101000010110";
rom_data(3253) <= "101000011000";
rom_data(3254) <= "101000011001";
rom_data(3255) <= "101000011011";
rom_data(3256) <= "101000011100";
rom_data(3257) <= "101000011110";
rom_data(3258) <= "101000100000";
rom_data(3259) <= "101000100001";
rom_data(3260) <= "101000100011";
rom_data(3261) <= "101000100100";
rom_data(3262) <= "101000100110";
rom_data(3263) <= "101000101000";
rom_data(3264) <= "101000101001";
rom_data(3265) <= "101000101011";
rom_data(3266) <= "101000101100";
rom_data(3267) <= "101000101110";
rom_data(3268) <= "101000110000";
rom_data(3269) <= "101000110001";
rom_data(3270) <= "101000110011";
rom_data(3271) <= "101000110100";
rom_data(3272) <= "101000110110";
rom_data(3273) <= "101000111000";
rom_data(3274) <= "101000111001";
rom_data(3275) <= "101000111011";
rom_data(3276) <= "101000111100";
rom_data(3277) <= "101000111110";
rom_data(3278) <= "101001000000";
rom_data(3279) <= "101001000001";
rom_data(3280) <= "101001000011";
rom_data(3281) <= "101001000100";
rom_data(3282) <= "101001000110";
rom_data(3283) <= "101001001000";
rom_data(3284) <= "101001001001";
rom_data(3285) <= "101001001011";
rom_data(3286) <= "101001001100";
rom_data(3287) <= "101001001110";
rom_data(3288) <= "101001010000";
rom_data(3289) <= "101001010001";
rom_data(3290) <= "101001010011";
rom_data(3291) <= "101001010100";
rom_data(3292) <= "101001010110";
rom_data(3293) <= "101001011000";
rom_data(3294) <= "101001011001";
rom_data(3295) <= "101001011011";
rom_data(3296) <= "101001011100";
rom_data(3297) <= "101001011110";
rom_data(3298) <= "101001100000";
rom_data(3299) <= "101001100001";
rom_data(3300) <= "101001100011";
rom_data(3301) <= "101001100100";
rom_data(3302) <= "101001100110";
rom_data(3303) <= "101001101000";
rom_data(3304) <= "101001101001";
rom_data(3305) <= "101001101011";
rom_data(3306) <= "101001101101";
rom_data(3307) <= "101001101110";
rom_data(3308) <= "101001110000";
rom_data(3309) <= "101001110001";
rom_data(3310) <= "101001110011";
rom_data(3311) <= "101001110101";
rom_data(3312) <= "101001110110";
rom_data(3313) <= "101001111000";
rom_data(3314) <= "101001111001";
rom_data(3315) <= "101001111011";
rom_data(3316) <= "101001111101";
rom_data(3317) <= "101001111110";
rom_data(3318) <= "101010000000";
rom_data(3319) <= "101010000010";
rom_data(3320) <= "101010000011";
rom_data(3321) <= "101010000101";
rom_data(3322) <= "101010000110";
rom_data(3323) <= "101010001000";
rom_data(3324) <= "101010001010";
rom_data(3325) <= "101010001011";
rom_data(3326) <= "101010001101";
rom_data(3327) <= "101010001111";
rom_data(3328) <= "101010010000";
rom_data(3329) <= "101010010010";
rom_data(3330) <= "101010010011";
rom_data(3331) <= "101010010101";
rom_data(3332) <= "101010010111";
rom_data(3333) <= "101010011000";
rom_data(3334) <= "101010011010";
rom_data(3335) <= "101010011100";
rom_data(3336) <= "101010011101";
rom_data(3337) <= "101010011111";
rom_data(3338) <= "101010100000";
rom_data(3339) <= "101010100010";
rom_data(3340) <= "101010100100";
rom_data(3341) <= "101010100101";
rom_data(3342) <= "101010100111";
rom_data(3343) <= "101010101001";
rom_data(3344) <= "101010101010";
rom_data(3345) <= "101010101100";
rom_data(3346) <= "101010101101";
rom_data(3347) <= "101010101111";
rom_data(3348) <= "101010110001";
rom_data(3349) <= "101010110010";
rom_data(3350) <= "101010110100";
rom_data(3351) <= "101010110110";
rom_data(3352) <= "101010110111";
rom_data(3353) <= "101010111001";
rom_data(3354) <= "101010111011";
rom_data(3355) <= "101010111100";
rom_data(3356) <= "101010111110";
rom_data(3357) <= "101011000000";
rom_data(3358) <= "101011000001";
rom_data(3359) <= "101011000011";
rom_data(3360) <= "101011000100";
rom_data(3361) <= "101011000110";
rom_data(3362) <= "101011001000";
rom_data(3363) <= "101011001001";
rom_data(3364) <= "101011001011";
rom_data(3365) <= "101011001101";
rom_data(3366) <= "101011001110";
rom_data(3367) <= "101011010000";
rom_data(3368) <= "101011010010";
rom_data(3369) <= "101011010011";
rom_data(3370) <= "101011010101";
rom_data(3371) <= "101011010111";
rom_data(3372) <= "101011011000";
rom_data(3373) <= "101011011010";
rom_data(3374) <= "101011011011";
rom_data(3375) <= "101011011101";
rom_data(3376) <= "101011011111";
rom_data(3377) <= "101011100000";
rom_data(3378) <= "101011100010";
rom_data(3379) <= "101011100100";
rom_data(3380) <= "101011100101";
rom_data(3381) <= "101011100111";
rom_data(3382) <= "101011101001";
rom_data(3383) <= "101011101010";
rom_data(3384) <= "101011101100";
rom_data(3385) <= "101011101110";
rom_data(3386) <= "101011101111";
rom_data(3387) <= "101011110001";
rom_data(3388) <= "101011110011";
rom_data(3389) <= "101011110100";
rom_data(3390) <= "101011110110";
rom_data(3391) <= "101011111000";
rom_data(3392) <= "101011111001";
rom_data(3393) <= "101011111011";
rom_data(3394) <= "101011111101";
rom_data(3395) <= "101011111110";
rom_data(3396) <= "101100000000";
rom_data(3397) <= "101100000001";
rom_data(3398) <= "101100000011";
rom_data(3399) <= "101100000101";
rom_data(3400) <= "101100000110";
rom_data(3401) <= "101100001000";
rom_data(3402) <= "101100001010";
rom_data(3403) <= "101100001011";
rom_data(3404) <= "101100001101";
rom_data(3405) <= "101100001111";
rom_data(3406) <= "101100010000";
rom_data(3407) <= "101100010010";
rom_data(3408) <= "101100010100";
rom_data(3409) <= "101100010101";
rom_data(3410) <= "101100010111";
rom_data(3411) <= "101100011001";
rom_data(3412) <= "101100011010";
rom_data(3413) <= "101100011100";
rom_data(3414) <= "101100011110";
rom_data(3415) <= "101100011111";
rom_data(3416) <= "101100100001";
rom_data(3417) <= "101100100011";
rom_data(3418) <= "101100100100";
rom_data(3419) <= "101100100110";
rom_data(3420) <= "101100101000";
rom_data(3421) <= "101100101001";
rom_data(3422) <= "101100101011";
rom_data(3423) <= "101100101101";
rom_data(3424) <= "101100101110";
rom_data(3425) <= "101100110000";
rom_data(3426) <= "101100110010";
rom_data(3427) <= "101100110011";
rom_data(3428) <= "101100110101";
rom_data(3429) <= "101100110111";
rom_data(3430) <= "101100111000";
rom_data(3431) <= "101100111010";
rom_data(3432) <= "101100111100";
rom_data(3433) <= "101100111110";
rom_data(3434) <= "101100111111";
rom_data(3435) <= "101101000001";
rom_data(3436) <= "101101000011";
rom_data(3437) <= "101101000100";
rom_data(3438) <= "101101000110";
rom_data(3439) <= "101101001000";
rom_data(3440) <= "101101001001";
rom_data(3441) <= "101101001011";
rom_data(3442) <= "101101001101";
rom_data(3443) <= "101101001110";
rom_data(3444) <= "101101010000";
rom_data(3445) <= "101101010010";
rom_data(3446) <= "101101010011";
rom_data(3447) <= "101101010101";
rom_data(3448) <= "101101010111";
rom_data(3449) <= "101101011000";
rom_data(3450) <= "101101011010";
rom_data(3451) <= "101101011100";
rom_data(3452) <= "101101011101";
rom_data(3453) <= "101101011111";
rom_data(3454) <= "101101100001";
rom_data(3455) <= "101101100011";
rom_data(3456) <= "101101100100";
rom_data(3457) <= "101101100110";
rom_data(3458) <= "101101101000";
rom_data(3459) <= "101101101001";
rom_data(3460) <= "101101101011";
rom_data(3461) <= "101101101101";
rom_data(3462) <= "101101101110";
rom_data(3463) <= "101101110000";
rom_data(3464) <= "101101110010";
rom_data(3465) <= "101101110011";
rom_data(3466) <= "101101110101";
rom_data(3467) <= "101101110111";
rom_data(3468) <= "101101111001";
rom_data(3469) <= "101101111010";
rom_data(3470) <= "101101111100";
rom_data(3471) <= "101101111110";
rom_data(3472) <= "101101111111";
rom_data(3473) <= "101110000001";
rom_data(3474) <= "101110000011";
rom_data(3475) <= "101110000100";
rom_data(3476) <= "101110000110";
rom_data(3477) <= "101110001000";
rom_data(3478) <= "101110001001";
rom_data(3479) <= "101110001011";
rom_data(3480) <= "101110001101";
rom_data(3481) <= "101110001111";
rom_data(3482) <= "101110010000";
rom_data(3483) <= "101110010010";
rom_data(3484) <= "101110010100";
rom_data(3485) <= "101110010101";
rom_data(3486) <= "101110010111";
rom_data(3487) <= "101110011001";
rom_data(3488) <= "101110011010";
rom_data(3489) <= "101110011100";
rom_data(3490) <= "101110011110";
rom_data(3491) <= "101110100000";
rom_data(3492) <= "101110100001";
rom_data(3493) <= "101110100011";
rom_data(3494) <= "101110100101";
rom_data(3495) <= "101110100110";
rom_data(3496) <= "101110101000";
rom_data(3497) <= "101110101010";
rom_data(3498) <= "101110101100";
rom_data(3499) <= "101110101101";
rom_data(3500) <= "101110101111";
rom_data(3501) <= "101110110001";
rom_data(3502) <= "101110110010";
rom_data(3503) <= "101110110100";
rom_data(3504) <= "101110110110";
rom_data(3505) <= "101110111000";
rom_data(3506) <= "101110111001";
rom_data(3507) <= "101110111011";
rom_data(3508) <= "101110111101";
rom_data(3509) <= "101110111110";
rom_data(3510) <= "101111000000";
rom_data(3511) <= "101111000010";
rom_data(3512) <= "101111000100";
rom_data(3513) <= "101111000101";
rom_data(3514) <= "101111000111";
rom_data(3515) <= "101111001001";
rom_data(3516) <= "101111001010";
rom_data(3517) <= "101111001100";
rom_data(3518) <= "101111001110";
rom_data(3519) <= "101111010000";
rom_data(3520) <= "101111010001";
rom_data(3521) <= "101111010011";
rom_data(3522) <= "101111010101";
rom_data(3523) <= "101111010110";
rom_data(3524) <= "101111011000";
rom_data(3525) <= "101111011010";
rom_data(3526) <= "101111011100";
rom_data(3527) <= "101111011101";
rom_data(3528) <= "101111011111";
rom_data(3529) <= "101111100001";
rom_data(3530) <= "101111100010";
rom_data(3531) <= "101111100100";
rom_data(3532) <= "101111100110";
rom_data(3533) <= "101111101000";
rom_data(3534) <= "101111101001";
rom_data(3535) <= "101111101011";
rom_data(3536) <= "101111101101";
rom_data(3537) <= "101111101111";
rom_data(3538) <= "101111110000";
rom_data(3539) <= "101111110010";
rom_data(3540) <= "101111110100";
rom_data(3541) <= "101111110101";
rom_data(3542) <= "101111110111";
rom_data(3543) <= "101111111001";
rom_data(3544) <= "101111111011";
rom_data(3545) <= "101111111100";
rom_data(3546) <= "101111111110";
rom_data(3547) <= "110000000000";
rom_data(3548) <= "110000000010";
rom_data(3549) <= "110000000011";
rom_data(3550) <= "110000000101";
rom_data(3551) <= "110000000111";
rom_data(3552) <= "110000001001";
rom_data(3553) <= "110000001010";
rom_data(3554) <= "110000001100";
rom_data(3555) <= "110000001110";
rom_data(3556) <= "110000001111";
rom_data(3557) <= "110000010001";
rom_data(3558) <= "110000010011";
rom_data(3559) <= "110000010101";
rom_data(3560) <= "110000010110";
rom_data(3561) <= "110000011000";
rom_data(3562) <= "110000011010";
rom_data(3563) <= "110000011100";
rom_data(3564) <= "110000011101";
rom_data(3565) <= "110000011111";
rom_data(3566) <= "110000100001";
rom_data(3567) <= "110000100011";
rom_data(3568) <= "110000100100";
rom_data(3569) <= "110000100110";
rom_data(3570) <= "110000101000";
rom_data(3571) <= "110000101010";
rom_data(3572) <= "110000101011";
rom_data(3573) <= "110000101101";
rom_data(3574) <= "110000101111";
rom_data(3575) <= "110000110001";
rom_data(3576) <= "110000110010";
rom_data(3577) <= "110000110100";
rom_data(3578) <= "110000110110";
rom_data(3579) <= "110000111000";
rom_data(3580) <= "110000111001";
rom_data(3581) <= "110000111011";
rom_data(3582) <= "110000111101";
rom_data(3583) <= "110000111111";
rom_data(3584) <= "110001000000";
rom_data(3585) <= "110001000010";
rom_data(3586) <= "110001000100";
rom_data(3587) <= "110001000110";
rom_data(3588) <= "110001000111";
rom_data(3589) <= "110001001001";
rom_data(3590) <= "110001001011";
rom_data(3591) <= "110001001101";
rom_data(3592) <= "110001001110";
rom_data(3593) <= "110001010000";
rom_data(3594) <= "110001010010";
rom_data(3595) <= "110001010100";
rom_data(3596) <= "110001010101";
rom_data(3597) <= "110001010111";
rom_data(3598) <= "110001011001";
rom_data(3599) <= "110001011011";
rom_data(3600) <= "110001011100";
rom_data(3601) <= "110001011110";
rom_data(3602) <= "110001100000";
rom_data(3603) <= "110001100010";
rom_data(3604) <= "110001100011";
rom_data(3605) <= "110001100101";
rom_data(3606) <= "110001100111";
rom_data(3607) <= "110001101001";
rom_data(3608) <= "110001101010";
rom_data(3609) <= "110001101100";
rom_data(3610) <= "110001101110";
rom_data(3611) <= "110001110000";
rom_data(3612) <= "110001110001";
rom_data(3613) <= "110001110011";
rom_data(3614) <= "110001110101";
rom_data(3615) <= "110001110111";
rom_data(3616) <= "110001111001";
rom_data(3617) <= "110001111010";
rom_data(3618) <= "110001111100";
rom_data(3619) <= "110001111110";
rom_data(3620) <= "110010000000";
rom_data(3621) <= "110010000001";
rom_data(3622) <= "110010000011";
rom_data(3623) <= "110010000101";
rom_data(3624) <= "110010000111";
rom_data(3625) <= "110010001000";
rom_data(3626) <= "110010001010";
rom_data(3627) <= "110010001100";
rom_data(3628) <= "110010001110";
rom_data(3629) <= "110010010000";
rom_data(3630) <= "110010010001";
rom_data(3631) <= "110010010011";
rom_data(3632) <= "110010010101";
rom_data(3633) <= "110010010111";
rom_data(3634) <= "110010011000";
rom_data(3635) <= "110010011010";
rom_data(3636) <= "110010011100";
rom_data(3637) <= "110010011110";
rom_data(3638) <= "110010100000";
rom_data(3639) <= "110010100001";
rom_data(3640) <= "110010100011";
rom_data(3641) <= "110010100101";
rom_data(3642) <= "110010100111";
rom_data(3643) <= "110010101000";
rom_data(3644) <= "110010101010";
rom_data(3645) <= "110010101100";
rom_data(3646) <= "110010101110";
rom_data(3647) <= "110010110000";
rom_data(3648) <= "110010110001";
rom_data(3649) <= "110010110011";
rom_data(3650) <= "110010110101";
rom_data(3651) <= "110010110111";
rom_data(3652) <= "110010111000";
rom_data(3653) <= "110010111010";
rom_data(3654) <= "110010111100";
rom_data(3655) <= "110010111110";
rom_data(3656) <= "110011000000";
rom_data(3657) <= "110011000001";
rom_data(3658) <= "110011000011";
rom_data(3659) <= "110011000101";
rom_data(3660) <= "110011000111";
rom_data(3661) <= "110011001000";
rom_data(3662) <= "110011001010";
rom_data(3663) <= "110011001100";
rom_data(3664) <= "110011001110";
rom_data(3665) <= "110011010000";
rom_data(3666) <= "110011010001";
rom_data(3667) <= "110011010011";
rom_data(3668) <= "110011010101";
rom_data(3669) <= "110011010111";
rom_data(3670) <= "110011011001";
rom_data(3671) <= "110011011010";
rom_data(3672) <= "110011011100";
rom_data(3673) <= "110011011110";
rom_data(3674) <= "110011100000";
rom_data(3675) <= "110011100010";
rom_data(3676) <= "110011100011";
rom_data(3677) <= "110011100101";
rom_data(3678) <= "110011100111";
rom_data(3679) <= "110011101001";
rom_data(3680) <= "110011101011";
rom_data(3681) <= "110011101100";
rom_data(3682) <= "110011101110";
rom_data(3683) <= "110011110000";
rom_data(3684) <= "110011110010";
rom_data(3685) <= "110011110100";
rom_data(3686) <= "110011110101";
rom_data(3687) <= "110011110111";
rom_data(3688) <= "110011111001";
rom_data(3689) <= "110011111011";
rom_data(3690) <= "110011111101";
rom_data(3691) <= "110011111110";
rom_data(3692) <= "110100000000";
rom_data(3693) <= "110100000010";
rom_data(3694) <= "110100000100";
rom_data(3695) <= "110100000110";
rom_data(3696) <= "110100000111";
rom_data(3697) <= "110100001001";
rom_data(3698) <= "110100001011";
rom_data(3699) <= "110100001101";
rom_data(3700) <= "110100001111";
rom_data(3701) <= "110100010000";
rom_data(3702) <= "110100010010";
rom_data(3703) <= "110100010100";
rom_data(3704) <= "110100010110";
rom_data(3705) <= "110100011000";
rom_data(3706) <= "110100011001";
rom_data(3707) <= "110100011011";
rom_data(3708) <= "110100011101";
rom_data(3709) <= "110100011111";
rom_data(3710) <= "110100100001";
rom_data(3711) <= "110100100011";
rom_data(3712) <= "110100100100";
rom_data(3713) <= "110100100110";
rom_data(3714) <= "110100101000";
rom_data(3715) <= "110100101010";
rom_data(3716) <= "110100101100";
rom_data(3717) <= "110100101101";
rom_data(3718) <= "110100101111";
rom_data(3719) <= "110100110001";
rom_data(3720) <= "110100110011";
rom_data(3721) <= "110100110101";
rom_data(3722) <= "110100110110";
rom_data(3723) <= "110100111000";
rom_data(3724) <= "110100111010";
rom_data(3725) <= "110100111100";
rom_data(3726) <= "110100111110";
rom_data(3727) <= "110101000000";
rom_data(3728) <= "110101000001";
rom_data(3729) <= "110101000011";
rom_data(3730) <= "110101000101";
rom_data(3731) <= "110101000111";
rom_data(3732) <= "110101001001";
rom_data(3733) <= "110101001011";
rom_data(3734) <= "110101001100";
rom_data(3735) <= "110101001110";
rom_data(3736) <= "110101010000";
rom_data(3737) <= "110101010010";
rom_data(3738) <= "110101010100";
rom_data(3739) <= "110101010101";
rom_data(3740) <= "110101010111";
rom_data(3741) <= "110101011001";
rom_data(3742) <= "110101011011";
rom_data(3743) <= "110101011101";
rom_data(3744) <= "110101011111";
rom_data(3745) <= "110101100000";
rom_data(3746) <= "110101100010";
rom_data(3747) <= "110101100100";
rom_data(3748) <= "110101100110";
rom_data(3749) <= "110101101000";
rom_data(3750) <= "110101101010";
rom_data(3751) <= "110101101011";
rom_data(3752) <= "110101101101";
rom_data(3753) <= "110101101111";
rom_data(3754) <= "110101110001";
rom_data(3755) <= "110101110011";
rom_data(3756) <= "110101110101";
rom_data(3757) <= "110101110110";
rom_data(3758) <= "110101111000";
rom_data(3759) <= "110101111010";
rom_data(3760) <= "110101111100";
rom_data(3761) <= "110101111110";
rom_data(3762) <= "110110000000";
rom_data(3763) <= "110110000001";
rom_data(3764) <= "110110000011";
rom_data(3765) <= "110110000101";
rom_data(3766) <= "110110000111";
rom_data(3767) <= "110110001001";
rom_data(3768) <= "110110001011";
rom_data(3769) <= "110110001100";
rom_data(3770) <= "110110001110";
rom_data(3771) <= "110110010000";
rom_data(3772) <= "110110010010";
rom_data(3773) <= "110110010100";
rom_data(3774) <= "110110010110";
rom_data(3775) <= "110110011000";
rom_data(3776) <= "110110011001";
rom_data(3777) <= "110110011011";
rom_data(3778) <= "110110011101";
rom_data(3779) <= "110110011111";
rom_data(3780) <= "110110100001";
rom_data(3781) <= "110110100011";
rom_data(3782) <= "110110100100";
rom_data(3783) <= "110110100110";
rom_data(3784) <= "110110101000";
rom_data(3785) <= "110110101010";
rom_data(3786) <= "110110101100";
rom_data(3787) <= "110110101110";
rom_data(3788) <= "110110110000";
rom_data(3789) <= "110110110001";
rom_data(3790) <= "110110110011";
rom_data(3791) <= "110110110101";
rom_data(3792) <= "110110110111";
rom_data(3793) <= "110110111001";
rom_data(3794) <= "110110111011";
rom_data(3795) <= "110110111100";
rom_data(3796) <= "110110111110";
rom_data(3797) <= "110111000000";
rom_data(3798) <= "110111000010";
rom_data(3799) <= "110111000100";
rom_data(3800) <= "110111000110";
rom_data(3801) <= "110111001000";
rom_data(3802) <= "110111001001";
rom_data(3803) <= "110111001011";
rom_data(3804) <= "110111001101";
rom_data(3805) <= "110111001111";
rom_data(3806) <= "110111010001";
rom_data(3807) <= "110111010011";
rom_data(3808) <= "110111010101";
rom_data(3809) <= "110111010110";
rom_data(3810) <= "110111011000";
rom_data(3811) <= "110111011010";
rom_data(3812) <= "110111011100";
rom_data(3813) <= "110111011110";
rom_data(3814) <= "110111100000";
rom_data(3815) <= "110111100010";
rom_data(3816) <= "110111100100";
rom_data(3817) <= "110111100101";
rom_data(3818) <= "110111100111";
rom_data(3819) <= "110111101001";
rom_data(3820) <= "110111101011";
rom_data(3821) <= "110111101101";
rom_data(3822) <= "110111101111";
rom_data(3823) <= "110111110001";
rom_data(3824) <= "110111110010";
rom_data(3825) <= "110111110100";
rom_data(3826) <= "110111110110";
rom_data(3827) <= "110111111000";
rom_data(3828) <= "110111111010";
rom_data(3829) <= "110111111100";
rom_data(3830) <= "110111111110";
rom_data(3831) <= "111000000000";
rom_data(3832) <= "111000000001";
rom_data(3833) <= "111000000011";
rom_data(3834) <= "111000000101";
rom_data(3835) <= "111000000111";
rom_data(3836) <= "111000001001";
rom_data(3837) <= "111000001011";
rom_data(3838) <= "111000001101";
rom_data(3839) <= "111000001111";
rom_data(3840) <= "111000010000";
rom_data(3841) <= "111000010010";
rom_data(3842) <= "111000010100";
rom_data(3843) <= "111000010110";
rom_data(3844) <= "111000011000";
rom_data(3845) <= "111000011010";
rom_data(3846) <= "111000011100";
rom_data(3847) <= "111000011110";
rom_data(3848) <= "111000011111";
rom_data(3849) <= "111000100001";
rom_data(3850) <= "111000100011";
rom_data(3851) <= "111000100101";
rom_data(3852) <= "111000100111";
rom_data(3853) <= "111000101001";
rom_data(3854) <= "111000101011";
rom_data(3855) <= "111000101101";
rom_data(3856) <= "111000101110";
rom_data(3857) <= "111000110000";
rom_data(3858) <= "111000110010";
rom_data(3859) <= "111000110100";
rom_data(3860) <= "111000110110";
rom_data(3861) <= "111000111000";
rom_data(3862) <= "111000111010";
rom_data(3863) <= "111000111100";
rom_data(3864) <= "111000111110";
rom_data(3865) <= "111000111111";
rom_data(3866) <= "111001000001";
rom_data(3867) <= "111001000011";
rom_data(3868) <= "111001000101";
rom_data(3869) <= "111001000111";
rom_data(3870) <= "111001001001";
rom_data(3871) <= "111001001011";
rom_data(3872) <= "111001001101";
rom_data(3873) <= "111001001111";
rom_data(3874) <= "111001010000";
rom_data(3875) <= "111001010010";
rom_data(3876) <= "111001010100";
rom_data(3877) <= "111001010110";
rom_data(3878) <= "111001011000";
rom_data(3879) <= "111001011010";
rom_data(3880) <= "111001011100";
rom_data(3881) <= "111001011110";
rom_data(3882) <= "111001100000";
rom_data(3883) <= "111001100001";
rom_data(3884) <= "111001100011";
rom_data(3885) <= "111001100101";
rom_data(3886) <= "111001100111";
rom_data(3887) <= "111001101001";
rom_data(3888) <= "111001101011";
rom_data(3889) <= "111001101101";
rom_data(3890) <= "111001101111";
rom_data(3891) <= "111001110001";
rom_data(3892) <= "111001110011";
rom_data(3893) <= "111001110100";
rom_data(3894) <= "111001110110";
rom_data(3895) <= "111001111000";
rom_data(3896) <= "111001111010";
rom_data(3897) <= "111001111100";
rom_data(3898) <= "111001111110";
rom_data(3899) <= "111010000000";
rom_data(3900) <= "111010000010";
rom_data(3901) <= "111010000100";
rom_data(3902) <= "111010000110";
rom_data(3903) <= "111010001000";
rom_data(3904) <= "111010001001";
rom_data(3905) <= "111010001011";
rom_data(3906) <= "111010001101";
rom_data(3907) <= "111010001111";
rom_data(3908) <= "111010010001";
rom_data(3909) <= "111010010011";
rom_data(3910) <= "111010010101";
rom_data(3911) <= "111010010111";
rom_data(3912) <= "111010011001";
rom_data(3913) <= "111010011011";
rom_data(3914) <= "111010011101";
rom_data(3915) <= "111010011110";
rom_data(3916) <= "111010100000";
rom_data(3917) <= "111010100010";
rom_data(3918) <= "111010100100";
rom_data(3919) <= "111010100110";
rom_data(3920) <= "111010101000";
rom_data(3921) <= "111010101010";
rom_data(3922) <= "111010101100";
rom_data(3923) <= "111010101110";
rom_data(3924) <= "111010110000";
rom_data(3925) <= "111010110010";
rom_data(3926) <= "111010110011";
rom_data(3927) <= "111010110101";
rom_data(3928) <= "111010110111";
rom_data(3929) <= "111010111001";
rom_data(3930) <= "111010111011";
rom_data(3931) <= "111010111101";
rom_data(3932) <= "111010111111";
rom_data(3933) <= "111011000001";
rom_data(3934) <= "111011000011";
rom_data(3935) <= "111011000101";
rom_data(3936) <= "111011000111";
rom_data(3937) <= "111011001001";
rom_data(3938) <= "111011001011";
rom_data(3939) <= "111011001100";
rom_data(3940) <= "111011001110";
rom_data(3941) <= "111011010000";
rom_data(3942) <= "111011010010";
rom_data(3943) <= "111011010100";
rom_data(3944) <= "111011010110";
rom_data(3945) <= "111011011000";
rom_data(3946) <= "111011011010";
rom_data(3947) <= "111011011100";
rom_data(3948) <= "111011011110";
rom_data(3949) <= "111011100000";
rom_data(3950) <= "111011100010";
rom_data(3951) <= "111011100100";
rom_data(3952) <= "111011100101";
rom_data(3953) <= "111011100111";
rom_data(3954) <= "111011101001";
rom_data(3955) <= "111011101011";
rom_data(3956) <= "111011101101";
rom_data(3957) <= "111011101111";
rom_data(3958) <= "111011110001";
rom_data(3959) <= "111011110011";
rom_data(3960) <= "111011110101";
rom_data(3961) <= "111011110111";
rom_data(3962) <= "111011111001";
rom_data(3963) <= "111011111011";
rom_data(3964) <= "111011111101";
rom_data(3965) <= "111011111111";
rom_data(3966) <= "111100000001";
rom_data(3967) <= "111100000011";
rom_data(3968) <= "111100000100";
rom_data(3969) <= "111100000110";
rom_data(3970) <= "111100001000";
rom_data(3971) <= "111100001010";
rom_data(3972) <= "111100001100";
rom_data(3973) <= "111100001110";
rom_data(3974) <= "111100010000";
rom_data(3975) <= "111100010010";
rom_data(3976) <= "111100010100";
rom_data(3977) <= "111100010110";
rom_data(3978) <= "111100011000";
rom_data(3979) <= "111100011010";
rom_data(3980) <= "111100011100";
rom_data(3981) <= "111100011110";
rom_data(3982) <= "111100100000";
rom_data(3983) <= "111100100010";
rom_data(3984) <= "111100100100";
rom_data(3985) <= "111100100101";
rom_data(3986) <= "111100100111";
rom_data(3987) <= "111100101001";
rom_data(3988) <= "111100101011";
rom_data(3989) <= "111100101101";
rom_data(3990) <= "111100101111";
rom_data(3991) <= "111100110001";
rom_data(3992) <= "111100110011";
rom_data(3993) <= "111100110101";
rom_data(3994) <= "111100110111";
rom_data(3995) <= "111100111001";
rom_data(3996) <= "111100111011";
rom_data(3997) <= "111100111101";
rom_data(3998) <= "111100111111";
rom_data(3999) <= "111101000001";
rom_data(4000) <= "111101000011";
rom_data(4001) <= "111101000101";
rom_data(4002) <= "111101000111";
rom_data(4003) <= "111101001001";
rom_data(4004) <= "111101001011";
rom_data(4005) <= "111101001100";
rom_data(4006) <= "111101001110";
rom_data(4007) <= "111101010000";
rom_data(4008) <= "111101010010";
rom_data(4009) <= "111101010100";
rom_data(4010) <= "111101010110";
rom_data(4011) <= "111101011000";
rom_data(4012) <= "111101011010";
rom_data(4013) <= "111101011100";
rom_data(4014) <= "111101011110";
rom_data(4015) <= "111101100000";
rom_data(4016) <= "111101100010";
rom_data(4017) <= "111101100100";
rom_data(4018) <= "111101100110";
rom_data(4019) <= "111101101000";
rom_data(4020) <= "111101101010";
rom_data(4021) <= "111101101100";
rom_data(4022) <= "111101101110";
rom_data(4023) <= "111101110000";
rom_data(4024) <= "111101110010";
rom_data(4025) <= "111101110100";
rom_data(4026) <= "111101110110";
rom_data(4027) <= "111101111000";
rom_data(4028) <= "111101111010";
rom_data(4029) <= "111101111100";
rom_data(4030) <= "111101111110";
rom_data(4031) <= "111110000000";
rom_data(4032) <= "111110000001";
rom_data(4033) <= "111110000011";
rom_data(4034) <= "111110000101";
rom_data(4035) <= "111110000111";
rom_data(4036) <= "111110001001";
rom_data(4037) <= "111110001011";
rom_data(4038) <= "111110001101";
rom_data(4039) <= "111110001111";
rom_data(4040) <= "111110010001";
rom_data(4041) <= "111110010011";
rom_data(4042) <= "111110010101";
rom_data(4043) <= "111110010111";
rom_data(4044) <= "111110011001";
rom_data(4045) <= "111110011011";
rom_data(4046) <= "111110011101";
rom_data(4047) <= "111110011111";
rom_data(4048) <= "111110100001";
rom_data(4049) <= "111110100011";
rom_data(4050) <= "111110100101";
rom_data(4051) <= "111110100111";
rom_data(4052) <= "111110101001";
rom_data(4053) <= "111110101011";
rom_data(4054) <= "111110101101";
rom_data(4055) <= "111110101111";
rom_data(4056) <= "111110110001";
rom_data(4057) <= "111110110011";
rom_data(4058) <= "111110110101";
rom_data(4059) <= "111110110111";
rom_data(4060) <= "111110111001";
rom_data(4061) <= "111110111011";
rom_data(4062) <= "111110111101";
rom_data(4063) <= "111110111111";
rom_data(4064) <= "111111000001";
rom_data(4065) <= "111111000011";
rom_data(4066) <= "111111000101";
rom_data(4067) <= "111111000111";
rom_data(4068) <= "111111001001";
rom_data(4069) <= "111111001011";
rom_data(4070) <= "111111001101";
rom_data(4071) <= "111111001111";
rom_data(4072) <= "111111010001";
rom_data(4073) <= "111111010011";
rom_data(4074) <= "111111010101";
rom_data(4075) <= "111111010111";
rom_data(4076) <= "111111011001";
rom_data(4077) <= "111111011011";
rom_data(4078) <= "111111011101";
rom_data(4079) <= "111111011111";
rom_data(4080) <= "111111100001";
rom_data(4081) <= "111111100011";
rom_data(4082) <= "111111100101";
rom_data(4083) <= "111111100111";
rom_data(4084) <= "111111101001";
rom_data(4085) <= "111111101011";
rom_data(4086) <= "111111101101";
rom_data(4087) <= "111111101111";
rom_data(4088) <= "111111110001";
rom_data(4089) <= "111111110011";
rom_data(4090) <= "111111110101";
rom_data(4091) <= "111111110111";
rom_data(4092) <= "111111111001";
rom_data(4093) <= "111111111011";
rom_data(4094) <= "111111111101";
rom_data(4095) <= "111111111111";


process(i_clk)
begin
	if rising_edge(i_clk) then
		if conv_integer(i_addr) < 4096 then
			o_data <= rom_data(conv_integer(i_addr));
		else
			o_data <= (others => '0');
		end if;
	end if;
end process;



end Behavioral;


