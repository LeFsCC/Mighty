library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;



entity rom_non_linear_mapper is
port ( 
	i_clk : in std_logic;
	i_addr : in std_logic_vector(9 downto 0);
	o_data : out std_logic_vector(11 downto 0)
);
end rom_non_linear_mapper;

architecture Behavioral of rom_non_linear_mapper is

TYPE ARRAY_ROM is array (natural range<>) of std_logic_vector(11 downto 0);

signal rom_data :ARRAY_ROM(1023 downto 0);

attribute RAM_STYLE : string;
attribute RAM_STYLE of rom_data: signal is "BLOCK";

begin


rom_data(0) <= "010100010111";
rom_data(1) <= "010100010111";
rom_data(2) <= "010100010111";
rom_data(3) <= "010100010111";
rom_data(4) <= "010100010111";
rom_data(5) <= "010100010111";
rom_data(6) <= "010100010111";
rom_data(7) <= "010100010111";
rom_data(8) <= "010100010111";
rom_data(9) <= "010100010111";
rom_data(10) <= "010100010111";
rom_data(11) <= "010100010111";
rom_data(12) <= "010100010111";
rom_data(13) <= "010100010111";
rom_data(14) <= "010100010111";
rom_data(15) <= "010100010111";
rom_data(16) <= "010100010111";
rom_data(17) <= "010100010111";
rom_data(18) <= "010100010111";
rom_data(19) <= "010100010111";
rom_data(20) <= "010100010111";
rom_data(21) <= "010100010111";
rom_data(22) <= "010100010111";
rom_data(23) <= "010100010111";
rom_data(24) <= "010100010111";
rom_data(25) <= "010100010111";
rom_data(26) <= "010100010111";
rom_data(27) <= "010100010111";
rom_data(28) <= "010100010111";
rom_data(29) <= "010100010111";
rom_data(30) <= "010100010111";
rom_data(31) <= "010100010111";
rom_data(32) <= "010100010111";
rom_data(33) <= "010100010111";
rom_data(34) <= "010100010111";
rom_data(35) <= "010100010111";
rom_data(36) <= "010100010111";
rom_data(37) <= "010100010111";
rom_data(38) <= "010100010111";
rom_data(39) <= "010100010111";
rom_data(40) <= "010100010111";
rom_data(41) <= "010100010111";
rom_data(42) <= "010100010111";
rom_data(43) <= "010100010111";
rom_data(44) <= "010100010111";
rom_data(45) <= "010100010111";
rom_data(46) <= "010100010111";
rom_data(47) <= "010100010111";
rom_data(48) <= "010100010111";
rom_data(49) <= "010100010111";
rom_data(50) <= "010100010111";
rom_data(51) <= "010100010111";
rom_data(52) <= "010100010111";
rom_data(53) <= "010100010111";
rom_data(54) <= "010100010111";
rom_data(55) <= "010100010111";
rom_data(56) <= "010100010111";
rom_data(57) <= "010100010111";
rom_data(58) <= "010100010111";
rom_data(59) <= "010100010111";
rom_data(60) <= "010100010111";
rom_data(61) <= "010100010111";
rom_data(62) <= "010100010111";
rom_data(63) <= "010100010111";
rom_data(64) <= "010100010111";
rom_data(65) <= "010100010111";
rom_data(66) <= "010100010111";
rom_data(67) <= "010100010111";
rom_data(68) <= "010100010111";
rom_data(69) <= "010100010111";
rom_data(70) <= "010100010111";
rom_data(71) <= "010100010111";
rom_data(72) <= "010100011000";
rom_data(73) <= "010100011000";
rom_data(74) <= "010100011000";
rom_data(75) <= "010100011000";
rom_data(76) <= "010100011000";
rom_data(77) <= "010100011000";
rom_data(78) <= "010100011000";
rom_data(79) <= "010100011000";
rom_data(80) <= "010100011000";
rom_data(81) <= "010100011000";
rom_data(82) <= "010100011000";
rom_data(83) <= "010100011000";
rom_data(84) <= "010100011000";
rom_data(85) <= "010100011000";
rom_data(86) <= "010100011000";
rom_data(87) <= "010100011000";
rom_data(88) <= "010100011000";
rom_data(89) <= "010100011000";
rom_data(90) <= "010100011000";
rom_data(91) <= "010100011000";
rom_data(92) <= "010100011000";
rom_data(93) <= "010100011000";
rom_data(94) <= "010100011000";
rom_data(95) <= "010100011000";
rom_data(96) <= "010100011000";
rom_data(97) <= "010100011000";
rom_data(98) <= "010100011000";
rom_data(99) <= "010100011000";
rom_data(100) <= "010100011000";
rom_data(101) <= "010100011000";
rom_data(102) <= "010100011001";
rom_data(103) <= "010100011001";
rom_data(104) <= "010100011001";
rom_data(105) <= "010100011001";
rom_data(106) <= "010100011001";
rom_data(107) <= "010100011001";
rom_data(108) <= "010100011001";
rom_data(109) <= "010100011001";
rom_data(110) <= "010100011001";
rom_data(111) <= "010100011001";
rom_data(112) <= "010100011001";
rom_data(113) <= "010100011001";
rom_data(114) <= "010100011001";
rom_data(115) <= "010100011001";
rom_data(116) <= "010100011001";
rom_data(117) <= "010100011001";
rom_data(118) <= "010100011001";
rom_data(119) <= "010100011001";
rom_data(120) <= "010100011001";
rom_data(121) <= "010100011001";
rom_data(122) <= "010100011001";
rom_data(123) <= "010100011001";
rom_data(124) <= "010100011001";
rom_data(125) <= "010100011010";
rom_data(126) <= "010100011010";
rom_data(127) <= "010100011010";
rom_data(128) <= "010100011010";
rom_data(129) <= "010100011010";
rom_data(130) <= "010100011010";
rom_data(131) <= "010100011010";
rom_data(132) <= "010100011010";
rom_data(133) <= "010100011010";
rom_data(134) <= "010100011010";
rom_data(135) <= "010100011010";
rom_data(136) <= "010100011010";
rom_data(137) <= "010100011010";
rom_data(138) <= "010100011010";
rom_data(139) <= "010100011010";
rom_data(140) <= "010100011010";
rom_data(141) <= "010100011010";
rom_data(142) <= "010100011010";
rom_data(143) <= "010100011010";
rom_data(144) <= "010100011011";
rom_data(145) <= "010100011011";
rom_data(146) <= "010100011011";
rom_data(147) <= "010100011011";
rom_data(148) <= "010100011011";
rom_data(149) <= "010100011011";
rom_data(150) <= "010100011011";
rom_data(151) <= "010100011011";
rom_data(152) <= "010100011011";
rom_data(153) <= "010100011011";
rom_data(154) <= "010100011011";
rom_data(155) <= "010100011011";
rom_data(156) <= "010100011011";
rom_data(157) <= "010100011011";
rom_data(158) <= "010100011011";
rom_data(159) <= "010100011011";
rom_data(160) <= "010100011011";
rom_data(161) <= "010100011100";
rom_data(162) <= "010100011100";
rom_data(163) <= "010100011100";
rom_data(164) <= "010100011100";
rom_data(165) <= "010100011100";
rom_data(166) <= "010100011100";
rom_data(167) <= "010100011100";
rom_data(168) <= "010100011100";
rom_data(169) <= "010100011100";
rom_data(170) <= "010100011100";
rom_data(171) <= "010100011100";
rom_data(172) <= "010100011100";
rom_data(173) <= "010100011100";
rom_data(174) <= "010100011100";
rom_data(175) <= "010100011100";
rom_data(176) <= "010100011100";
rom_data(177) <= "010100011101";
rom_data(178) <= "010100011101";
rom_data(179) <= "010100011101";
rom_data(180) <= "010100011101";
rom_data(181) <= "010100011101";
rom_data(182) <= "010100011101";
rom_data(183) <= "010100011101";
rom_data(184) <= "010100011101";
rom_data(185) <= "010100011101";
rom_data(186) <= "010100011101";
rom_data(187) <= "010100011101";
rom_data(188) <= "010100011101";
rom_data(189) <= "010100011101";
rom_data(190) <= "010100011101";
rom_data(191) <= "010100011110";
rom_data(192) <= "010100011110";
rom_data(193) <= "010100011110";
rom_data(194) <= "010100011110";
rom_data(195) <= "010100011110";
rom_data(196) <= "010100011110";
rom_data(197) <= "010100011110";
rom_data(198) <= "010100011110";
rom_data(199) <= "010100011110";
rom_data(200) <= "010100011110";
rom_data(201) <= "010100011110";
rom_data(202) <= "010100011110";
rom_data(203) <= "010100011110";
rom_data(204) <= "010100011111";
rom_data(205) <= "010100011111";
rom_data(206) <= "010100011111";
rom_data(207) <= "010100011111";
rom_data(208) <= "010100011111";
rom_data(209) <= "010100011111";
rom_data(210) <= "010100011111";
rom_data(211) <= "010100011111";
rom_data(212) <= "010100011111";
rom_data(213) <= "010100011111";
rom_data(214) <= "010100011111";
rom_data(215) <= "010100011111";
rom_data(216) <= "010100100000";
rom_data(217) <= "010100100000";
rom_data(218) <= "010100100000";
rom_data(219) <= "010100100000";
rom_data(220) <= "010100100000";
rom_data(221) <= "010100100000";
rom_data(222) <= "010100100000";
rom_data(223) <= "010100100000";
rom_data(224) <= "010100100000";
rom_data(225) <= "010100100000";
rom_data(226) <= "010100100000";
rom_data(227) <= "010100100000";
rom_data(228) <= "010100100001";
rom_data(229) <= "010100100001";
rom_data(230) <= "010100100001";
rom_data(231) <= "010100100001";
rom_data(232) <= "010100100001";
rom_data(233) <= "010100100001";
rom_data(234) <= "010100100001";
rom_data(235) <= "010100100001";
rom_data(236) <= "010100100001";
rom_data(237) <= "010100100001";
rom_data(238) <= "010100100001";
rom_data(239) <= "010100100010";
rom_data(240) <= "010100100010";
rom_data(241) <= "010100100010";
rom_data(242) <= "010100100010";
rom_data(243) <= "010100100010";
rom_data(244) <= "010100100010";
rom_data(245) <= "010100100010";
rom_data(246) <= "010100100010";
rom_data(247) <= "010100100010";
rom_data(248) <= "010100100010";
rom_data(249) <= "010100100010";
rom_data(250) <= "010100100011";
rom_data(251) <= "010100100011";
rom_data(252) <= "010100100011";
rom_data(253) <= "010100100011";
rom_data(254) <= "010100100011";
rom_data(255) <= "010100100011";
rom_data(256) <= "010100100011";
rom_data(257) <= "010100100011";
rom_data(258) <= "010100100011";
rom_data(259) <= "010100100011";
rom_data(260) <= "010100100100";
rom_data(261) <= "010100100100";
rom_data(262) <= "010100100100";
rom_data(263) <= "010100100100";
rom_data(264) <= "010100100100";
rom_data(265) <= "010100100100";
rom_data(266) <= "010100100100";
rom_data(267) <= "010100100100";
rom_data(268) <= "010100100100";
rom_data(269) <= "010100100100";
rom_data(270) <= "010100100101";
rom_data(271) <= "010100100101";
rom_data(272) <= "010100100101";
rom_data(273) <= "010100100101";
rom_data(274) <= "010100100101";
rom_data(275) <= "010100100101";
rom_data(276) <= "010100100101";
rom_data(277) <= "010100100101";
rom_data(278) <= "010100100101";
rom_data(279) <= "010100100110";
rom_data(280) <= "010100100110";
rom_data(281) <= "010100100110";
rom_data(282) <= "010100100110";
rom_data(283) <= "010100100110";
rom_data(284) <= "010100100110";
rom_data(285) <= "010100100110";
rom_data(286) <= "010100100110";
rom_data(287) <= "010100100110";
rom_data(288) <= "010100100111";
rom_data(289) <= "010100100111";
rom_data(290) <= "010100100111";
rom_data(291) <= "010100100111";
rom_data(292) <= "010100100111";
rom_data(293) <= "010100100111";
rom_data(294) <= "010100100111";
rom_data(295) <= "010100100111";
rom_data(296) <= "010100100111";
rom_data(297) <= "010100101000";
rom_data(298) <= "010100101000";
rom_data(299) <= "010100101000";
rom_data(300) <= "010100101000";
rom_data(301) <= "010100101000";
rom_data(302) <= "010100101000";
rom_data(303) <= "010100101000";
rom_data(304) <= "010100101000";
rom_data(305) <= "010100101000";
rom_data(306) <= "010100101001";
rom_data(307) <= "010100101001";
rom_data(308) <= "010100101001";
rom_data(309) <= "010100101001";
rom_data(310) <= "010100101001";
rom_data(311) <= "010100101001";
rom_data(312) <= "010100101001";
rom_data(313) <= "010100101001";
rom_data(314) <= "010100101010";
rom_data(315) <= "010100101010";
rom_data(316) <= "010100101010";
rom_data(317) <= "010100101010";
rom_data(318) <= "010100101010";
rom_data(319) <= "010100101010";
rom_data(320) <= "010100101010";
rom_data(321) <= "010100101010";
rom_data(322) <= "010100101011";
rom_data(323) <= "010100101011";
rom_data(324) <= "010100101011";
rom_data(325) <= "010100101011";
rom_data(326) <= "010100101011";
rom_data(327) <= "010100101011";
rom_data(328) <= "010100101011";
rom_data(329) <= "010100101011";
rom_data(330) <= "010100101100";
rom_data(331) <= "010100101100";
rom_data(332) <= "010100101100";
rom_data(333) <= "010100101100";
rom_data(334) <= "010100101100";
rom_data(335) <= "010100101100";
rom_data(336) <= "010100101100";
rom_data(337) <= "010100101100";
rom_data(338) <= "010100101101";
rom_data(339) <= "010100101101";
rom_data(340) <= "010100101101";
rom_data(341) <= "010100101101";
rom_data(342) <= "010100101101";
rom_data(343) <= "010100101101";
rom_data(344) <= "010100101101";
rom_data(345) <= "010100101101";
rom_data(346) <= "010100101110";
rom_data(347) <= "010100101110";
rom_data(348) <= "010100101110";
rom_data(349) <= "010100101110";
rom_data(350) <= "010100101110";
rom_data(351) <= "010100101110";
rom_data(352) <= "010100101110";
rom_data(353) <= "010100101111";
rom_data(354) <= "010100101111";
rom_data(355) <= "010100101111";
rom_data(356) <= "010100101111";
rom_data(357) <= "010100101111";
rom_data(358) <= "010100101111";
rom_data(359) <= "010100101111";
rom_data(360) <= "010100110000";
rom_data(361) <= "010100110000";
rom_data(362) <= "010100110000";
rom_data(363) <= "010100110000";
rom_data(364) <= "010100110000";
rom_data(365) <= "010100110000";
rom_data(366) <= "010100110000";
rom_data(367) <= "010100110000";
rom_data(368) <= "010100110001";
rom_data(369) <= "010100110001";
rom_data(370) <= "010100110001";
rom_data(371) <= "010100110001";
rom_data(372) <= "010100110001";
rom_data(373) <= "010100110001";
rom_data(374) <= "010100110001";
rom_data(375) <= "010100110010";
rom_data(376) <= "010100110010";
rom_data(377) <= "010100110010";
rom_data(378) <= "010100110010";
rom_data(379) <= "010100110010";
rom_data(380) <= "010100110010";
rom_data(381) <= "010100110011";
rom_data(382) <= "010100110011";
rom_data(383) <= "010100110011";
rom_data(384) <= "010100110011";
rom_data(385) <= "010100110011";
rom_data(386) <= "010100110011";
rom_data(387) <= "010100110011";
rom_data(388) <= "010100110100";
rom_data(389) <= "010100110100";
rom_data(390) <= "010100110100";
rom_data(391) <= "010100110100";
rom_data(392) <= "010100110100";
rom_data(393) <= "010100110100";
rom_data(394) <= "010100110100";
rom_data(395) <= "010100110101";
rom_data(396) <= "010100110101";
rom_data(397) <= "010100110101";
rom_data(398) <= "010100110101";
rom_data(399) <= "010100110101";
rom_data(400) <= "010100110101";
rom_data(401) <= "010100110110";
rom_data(402) <= "010100110110";
rom_data(403) <= "010100110110";
rom_data(404) <= "010100110110";
rom_data(405) <= "010100110110";
rom_data(406) <= "010100110110";
rom_data(407) <= "010100110110";
rom_data(408) <= "010100110111";
rom_data(409) <= "010100110111";
rom_data(410) <= "010100110111";
rom_data(411) <= "010100110111";
rom_data(412) <= "010100110111";
rom_data(413) <= "010100110111";
rom_data(414) <= "010100111000";
rom_data(415) <= "010100111000";
rom_data(416) <= "010100111000";
rom_data(417) <= "010100111000";
rom_data(418) <= "010100111000";
rom_data(419) <= "010100111000";
rom_data(420) <= "010100111001";
rom_data(421) <= "010100111001";
rom_data(422) <= "010100111001";
rom_data(423) <= "010100111001";
rom_data(424) <= "010100111001";
rom_data(425) <= "010100111001";
rom_data(426) <= "010100111010";
rom_data(427) <= "010100111010";
rom_data(428) <= "010100111010";
rom_data(429) <= "010100111010";
rom_data(430) <= "010100111010";
rom_data(431) <= "010100111010";
rom_data(432) <= "010100111011";
rom_data(433) <= "010100111011";
rom_data(434) <= "010100111011";
rom_data(435) <= "010100111011";
rom_data(436) <= "010100111011";
rom_data(437) <= "010100111011";
rom_data(438) <= "010100111100";
rom_data(439) <= "010100111100";
rom_data(440) <= "010100111100";
rom_data(441) <= "010100111100";
rom_data(442) <= "010100111100";
rom_data(443) <= "010100111100";
rom_data(444) <= "010100111101";
rom_data(445) <= "010100111101";
rom_data(446) <= "010100111101";
rom_data(447) <= "010100111101";
rom_data(448) <= "010100111101";
rom_data(449) <= "010100111101";
rom_data(450) <= "010100111110";
rom_data(451) <= "010100111110";
rom_data(452) <= "010100111110";
rom_data(453) <= "010100111110";
rom_data(454) <= "010100111110";
rom_data(455) <= "010100111110";
rom_data(456) <= "010100111111";
rom_data(457) <= "010100111111";
rom_data(458) <= "010100111111";
rom_data(459) <= "010100111111";
rom_data(460) <= "010100111111";
rom_data(461) <= "010101000000";
rom_data(462) <= "010101000000";
rom_data(463) <= "010101000000";
rom_data(464) <= "010101000000";
rom_data(465) <= "010101000000";
rom_data(466) <= "010101000000";
rom_data(467) <= "010101000001";
rom_data(468) <= "010101000001";
rom_data(469) <= "010101000001";
rom_data(470) <= "010101000001";
rom_data(471) <= "010101000001";
rom_data(472) <= "010101000010";
rom_data(473) <= "010101000010";
rom_data(474) <= "010101000010";
rom_data(475) <= "010101000010";
rom_data(476) <= "010101000010";
rom_data(477) <= "010101000010";
rom_data(478) <= "010101000011";
rom_data(479) <= "010101000011";
rom_data(480) <= "010101000011";
rom_data(481) <= "010101000011";
rom_data(482) <= "010101000011";
rom_data(483) <= "010101000100";
rom_data(484) <= "010101000100";
rom_data(485) <= "010101000100";
rom_data(486) <= "010101000100";
rom_data(487) <= "010101000100";
rom_data(488) <= "010101000100";
rom_data(489) <= "010101000101";
rom_data(490) <= "010101000101";
rom_data(491) <= "010101000101";
rom_data(492) <= "010101000101";
rom_data(493) <= "010101000101";
rom_data(494) <= "010101000110";
rom_data(495) <= "010101000110";
rom_data(496) <= "010101000110";
rom_data(497) <= "010101000110";
rom_data(498) <= "010101000110";
rom_data(499) <= "010101000111";
rom_data(500) <= "010101000111";
rom_data(501) <= "010101000111";
rom_data(502) <= "010101000111";
rom_data(503) <= "010101000111";
rom_data(504) <= "010101001000";
rom_data(505) <= "010101001000";
rom_data(506) <= "010101001000";
rom_data(507) <= "010101001000";
rom_data(508) <= "010101001000";
rom_data(509) <= "010101001001";
rom_data(510) <= "010101001001";
rom_data(511) <= "010101001001";
rom_data(512) <= "010101001001";
rom_data(513) <= "010101001001";
rom_data(514) <= "010101001001";
rom_data(515) <= "010101001010";
rom_data(516) <= "010101001010";
rom_data(517) <= "010101001010";
rom_data(518) <= "010101001010";
rom_data(519) <= "010101001010";
rom_data(520) <= "010101001011";
rom_data(521) <= "010101001011";
rom_data(522) <= "010101001011";
rom_data(523) <= "010101001011";
rom_data(524) <= "010101001011";
rom_data(525) <= "010101001100";
rom_data(526) <= "010101001100";
rom_data(527) <= "010101001100";
rom_data(528) <= "010101001100";
rom_data(529) <= "010101001101";
rom_data(530) <= "010101001101";
rom_data(531) <= "010101001101";
rom_data(532) <= "010101001101";
rom_data(533) <= "010101001101";
rom_data(534) <= "010101001110";
rom_data(535) <= "010101001110";
rom_data(536) <= "010101001110";
rom_data(537) <= "010101001110";
rom_data(538) <= "010101001110";
rom_data(539) <= "010101001111";
rom_data(540) <= "010101001111";
rom_data(541) <= "010101001111";
rom_data(542) <= "010101001111";
rom_data(543) <= "010101001111";
rom_data(544) <= "010101010000";
rom_data(545) <= "010101010000";
rom_data(546) <= "010101010000";
rom_data(547) <= "010101010000";
rom_data(548) <= "010101010000";
rom_data(549) <= "010101010001";
rom_data(550) <= "010101010001";
rom_data(551) <= "010101010001";
rom_data(552) <= "010101010001";
rom_data(553) <= "010101010010";
rom_data(554) <= "010101010010";
rom_data(555) <= "010101010010";
rom_data(556) <= "010101010010";
rom_data(557) <= "010101010010";
rom_data(558) <= "010101010011";
rom_data(559) <= "010101010011";
rom_data(560) <= "010101010011";
rom_data(561) <= "010101010011";
rom_data(562) <= "010101010011";
rom_data(563) <= "010101010100";
rom_data(564) <= "010101010100";
rom_data(565) <= "010101010100";
rom_data(566) <= "010101010100";
rom_data(567) <= "010101010101";
rom_data(568) <= "010101010101";
rom_data(569) <= "010101010101";
rom_data(570) <= "010101010101";
rom_data(571) <= "010101010101";
rom_data(572) <= "010101010110";
rom_data(573) <= "010101010110";
rom_data(574) <= "010101010110";
rom_data(575) <= "010101010110";
rom_data(576) <= "010101010111";
rom_data(577) <= "010101010111";
rom_data(578) <= "010101010111";
rom_data(579) <= "010101010111";
rom_data(580) <= "010101010111";
rom_data(581) <= "010101011000";
rom_data(582) <= "010101011000";
rom_data(583) <= "010101011000";
rom_data(584) <= "010101011000";
rom_data(585) <= "010101011001";
rom_data(586) <= "010101011001";
rom_data(587) <= "010101011001";
rom_data(588) <= "010101011001";
rom_data(589) <= "010101011001";
rom_data(590) <= "010101011010";
rom_data(591) <= "010101011010";
rom_data(592) <= "010101011010";
rom_data(593) <= "010101011010";
rom_data(594) <= "010101011011";
rom_data(595) <= "010101011011";
rom_data(596) <= "010101011011";
rom_data(597) <= "010101011011";
rom_data(598) <= "010101011100";
rom_data(599) <= "010101011100";
rom_data(600) <= "010101011100";
rom_data(601) <= "010101011100";
rom_data(602) <= "010101011100";
rom_data(603) <= "010101011101";
rom_data(604) <= "010101011101";
rom_data(605) <= "010101011101";
rom_data(606) <= "010101011101";
rom_data(607) <= "010101011110";
rom_data(608) <= "010101011110";
rom_data(609) <= "010101011110";
rom_data(610) <= "010101011110";
rom_data(611) <= "010101011111";
rom_data(612) <= "010101011111";
rom_data(613) <= "010101011111";
rom_data(614) <= "010101011111";
rom_data(615) <= "010101100000";
rom_data(616) <= "010101100000";
rom_data(617) <= "010101100000";
rom_data(618) <= "010101100000";
rom_data(619) <= "010101100000";
rom_data(620) <= "010101100001";
rom_data(621) <= "010101100001";
rom_data(622) <= "010101100001";
rom_data(623) <= "010101100001";
rom_data(624) <= "010101100010";
rom_data(625) <= "010101100010";
rom_data(626) <= "010101100010";
rom_data(627) <= "010101100010";
rom_data(628) <= "010101100011";
rom_data(629) <= "010101100011";
rom_data(630) <= "010101100011";
rom_data(631) <= "010101100011";
rom_data(632) <= "010101100100";
rom_data(633) <= "010101100100";
rom_data(634) <= "010101100100";
rom_data(635) <= "010101100100";
rom_data(636) <= "010101100101";
rom_data(637) <= "010101100101";
rom_data(638) <= "010101100101";
rom_data(639) <= "010101100101";
rom_data(640) <= "010101100110";
rom_data(641) <= "010101100110";
rom_data(642) <= "010101100110";
rom_data(643) <= "010101100110";
rom_data(644) <= "010101100111";
rom_data(645) <= "010101100111";
rom_data(646) <= "010101100111";
rom_data(647) <= "010101100111";
rom_data(648) <= "010101101000";
rom_data(649) <= "010101101000";
rom_data(650) <= "010101101000";
rom_data(651) <= "010101101000";
rom_data(652) <= "010101101001";
rom_data(653) <= "010101101001";
rom_data(654) <= "010101101001";
rom_data(655) <= "010101101001";
rom_data(656) <= "010101101010";
rom_data(657) <= "010101101010";
rom_data(658) <= "010101101010";
rom_data(659) <= "010101101010";
rom_data(660) <= "010101101011";
rom_data(661) <= "010101101011";
rom_data(662) <= "010101101011";
rom_data(663) <= "010101101011";
rom_data(664) <= "010101101100";
rom_data(665) <= "010101101100";
rom_data(666) <= "010101101100";
rom_data(667) <= "010101101100";
rom_data(668) <= "010101101101";
rom_data(669) <= "010101101101";
rom_data(670) <= "010101101101";
rom_data(671) <= "010101101101";
rom_data(672) <= "010101101110";
rom_data(673) <= "010101101110";
rom_data(674) <= "010101101110";
rom_data(675) <= "010101101110";
rom_data(676) <= "010101101111";
rom_data(677) <= "010101101111";
rom_data(678) <= "010101101111";
rom_data(679) <= "010101101111";
rom_data(680) <= "010101110000";
rom_data(681) <= "010101110000";
rom_data(682) <= "010101110000";
rom_data(683) <= "010101110001";
rom_data(684) <= "010101110001";
rom_data(685) <= "010101110001";
rom_data(686) <= "010101110001";
rom_data(687) <= "010101110010";
rom_data(688) <= "010101110010";
rom_data(689) <= "010101110010";
rom_data(690) <= "010101110010";
rom_data(691) <= "010101110011";
rom_data(692) <= "010101110011";
rom_data(693) <= "010101110011";
rom_data(694) <= "010101110011";
rom_data(695) <= "010101110100";
rom_data(696) <= "010101110100";
rom_data(697) <= "010101110100";
rom_data(698) <= "010101110101";
rom_data(699) <= "010101110101";
rom_data(700) <= "010101110101";
rom_data(701) <= "010101110101";
rom_data(702) <= "010101110110";
rom_data(703) <= "010101110110";
rom_data(704) <= "010101110110";
rom_data(705) <= "010101110110";
rom_data(706) <= "010101110111";
rom_data(707) <= "010101110111";
rom_data(708) <= "010101110111";
rom_data(709) <= "010101111000";
rom_data(710) <= "010101111000";
rom_data(711) <= "010101111000";
rom_data(712) <= "010101111000";
rom_data(713) <= "010101111001";
rom_data(714) <= "010101111001";
rom_data(715) <= "010101111001";
rom_data(716) <= "010101111001";
rom_data(717) <= "010101111010";
rom_data(718) <= "010101111010";
rom_data(719) <= "010101111010";
rom_data(720) <= "010101111011";
rom_data(721) <= "010101111011";
rom_data(722) <= "010101111011";
rom_data(723) <= "010101111011";
rom_data(724) <= "010101111100";
rom_data(725) <= "010101111100";
rom_data(726) <= "010101111100";
rom_data(727) <= "010101111101";
rom_data(728) <= "010101111101";
rom_data(729) <= "010101111101";
rom_data(730) <= "010101111101";
rom_data(731) <= "010101111110";
rom_data(732) <= "010101111110";
rom_data(733) <= "010101111110";
rom_data(734) <= "010101111110";
rom_data(735) <= "010101111111";
rom_data(736) <= "010101111111";
rom_data(737) <= "010101111111";
rom_data(738) <= "010110000000";
rom_data(739) <= "010110000000";
rom_data(740) <= "010110000000";
rom_data(741) <= "010110000000";
rom_data(742) <= "010110000001";
rom_data(743) <= "010110000001";
rom_data(744) <= "010110000001";
rom_data(745) <= "010110000010";
rom_data(746) <= "010110000010";
rom_data(747) <= "010110000010";
rom_data(748) <= "010110000010";
rom_data(749) <= "010110000011";
rom_data(750) <= "010110000011";
rom_data(751) <= "010110000011";
rom_data(752) <= "010110000100";
rom_data(753) <= "010110000100";
rom_data(754) <= "010110000100";
rom_data(755) <= "010110000101";
rom_data(756) <= "010110000101";
rom_data(757) <= "010110000101";
rom_data(758) <= "010110000101";
rom_data(759) <= "010110000110";
rom_data(760) <= "010110000110";
rom_data(761) <= "010110000110";
rom_data(762) <= "010110000111";
rom_data(763) <= "010110000111";
rom_data(764) <= "010110000111";
rom_data(765) <= "010110000111";
rom_data(766) <= "010110001000";
rom_data(767) <= "010110001000";
rom_data(768) <= "010110001000";
rom_data(769) <= "010110001001";
rom_data(770) <= "010110001001";
rom_data(771) <= "010110001001";
rom_data(772) <= "010110001010";
rom_data(773) <= "010110001010";
rom_data(774) <= "010110001010";
rom_data(775) <= "010110001010";
rom_data(776) <= "010110001011";
rom_data(777) <= "010110001011";
rom_data(778) <= "010110001011";
rom_data(779) <= "010110001100";
rom_data(780) <= "010110001100";
rom_data(781) <= "010110001100";
rom_data(782) <= "010110001101";
rom_data(783) <= "010110001101";
rom_data(784) <= "010110001101";
rom_data(785) <= "010110001101";
rom_data(786) <= "010110001110";
rom_data(787) <= "010110001110";
rom_data(788) <= "010110001110";
rom_data(789) <= "010110001111";
rom_data(790) <= "010110001111";
rom_data(791) <= "010110001111";
rom_data(792) <= "010110010000";
rom_data(793) <= "010110010000";
rom_data(794) <= "010110010000";
rom_data(795) <= "010110010000";
rom_data(796) <= "010110010001";
rom_data(797) <= "010110010001";
rom_data(798) <= "010110010001";
rom_data(799) <= "010110010010";
rom_data(800) <= "010110010010";
rom_data(801) <= "010110010010";
rom_data(802) <= "010110010011";
rom_data(803) <= "010110010011";
rom_data(804) <= "010110010011";
rom_data(805) <= "010110010100";
rom_data(806) <= "010110010100";
rom_data(807) <= "010110010100";
rom_data(808) <= "010110010101";
rom_data(809) <= "010110010101";
rom_data(810) <= "010110010101";
rom_data(811) <= "010110010101";
rom_data(812) <= "010110010110";
rom_data(813) <= "010110010110";
rom_data(814) <= "010110010110";
rom_data(815) <= "010110010111";
rom_data(816) <= "010110010111";
rom_data(817) <= "010110010111";
rom_data(818) <= "010110011000";
rom_data(819) <= "010110011000";
rom_data(820) <= "010110011000";
rom_data(821) <= "010110011001";
rom_data(822) <= "010110011001";
rom_data(823) <= "010110011001";
rom_data(824) <= "010110011010";
rom_data(825) <= "010110011010";
rom_data(826) <= "010110011010";
rom_data(827) <= "010110011011";
rom_data(828) <= "010110011011";
rom_data(829) <= "010110011011";
rom_data(830) <= "010110011011";
rom_data(831) <= "010110011100";
rom_data(832) <= "010110011100";
rom_data(833) <= "010110011100";
rom_data(834) <= "010110011101";
rom_data(835) <= "010110011101";
rom_data(836) <= "010110011101";
rom_data(837) <= "010110011110";
rom_data(838) <= "010110011110";
rom_data(839) <= "010110011110";
rom_data(840) <= "010110011111";
rom_data(841) <= "010110011111";
rom_data(842) <= "010110011111";
rom_data(843) <= "010110100000";
rom_data(844) <= "010110100000";
rom_data(845) <= "010110100000";
rom_data(846) <= "010110100001";
rom_data(847) <= "010110100001";
rom_data(848) <= "010110100001";
rom_data(849) <= "010110100010";
rom_data(850) <= "010110100010";
rom_data(851) <= "010110100010";
rom_data(852) <= "010110100011";
rom_data(853) <= "010110100011";
rom_data(854) <= "010110100011";
rom_data(855) <= "010110100100";
rom_data(856) <= "010110100100";
rom_data(857) <= "010110100100";
rom_data(858) <= "010110100101";
rom_data(859) <= "010110100101";
rom_data(860) <= "010110100101";
rom_data(861) <= "010110100110";
rom_data(862) <= "010110100110";
rom_data(863) <= "010110100110";
rom_data(864) <= "010110100111";
rom_data(865) <= "010110100111";
rom_data(866) <= "010110100111";
rom_data(867) <= "010110101000";
rom_data(868) <= "010110101000";
rom_data(869) <= "010110101000";
rom_data(870) <= "010110101001";
rom_data(871) <= "010110101001";
rom_data(872) <= "010110101001";
rom_data(873) <= "010110101010";
rom_data(874) <= "010110101010";
rom_data(875) <= "010110101010";
rom_data(876) <= "010110101011";
rom_data(877) <= "010110101011";
rom_data(878) <= "010110101011";
rom_data(879) <= "010110101100";
rom_data(880) <= "010110101100";
rom_data(881) <= "010110101100";
rom_data(882) <= "010110101101";
rom_data(883) <= "010110101101";
rom_data(884) <= "010110101101";
rom_data(885) <= "010110101110";
rom_data(886) <= "010110101110";
rom_data(887) <= "010110101110";
rom_data(888) <= "010110101111";
rom_data(889) <= "010110101111";
rom_data(890) <= "010110101111";
rom_data(891) <= "010110110000";
rom_data(892) <= "010110110000";
rom_data(893) <= "010110110000";
rom_data(894) <= "010110110001";
rom_data(895) <= "010110110001";
rom_data(896) <= "010110110001";
rom_data(897) <= "010110110010";
rom_data(898) <= "010110110010";
rom_data(899) <= "010110110010";
rom_data(900) <= "010110110011";
rom_data(901) <= "010110110011";
rom_data(902) <= "010110110100";
rom_data(903) <= "010110110100";
rom_data(904) <= "010110110100";
rom_data(905) <= "010110110101";
rom_data(906) <= "010110110101";
rom_data(907) <= "010110110101";
rom_data(908) <= "010110110110";
rom_data(909) <= "010110110110";
rom_data(910) <= "010110110110";
rom_data(911) <= "010110110111";
rom_data(912) <= "010110110111";
rom_data(913) <= "010110110111";
rom_data(914) <= "010110111000";
rom_data(915) <= "010110111000";
rom_data(916) <= "010110111000";
rom_data(917) <= "010110111001";
rom_data(918) <= "010110111001";
rom_data(919) <= "010110111010";
rom_data(920) <= "010110111010";
rom_data(921) <= "010110111010";
rom_data(922) <= "010110111011";
rom_data(923) <= "010110111011";
rom_data(924) <= "010110111011";
rom_data(925) <= "010110111100";
rom_data(926) <= "010110111100";
rom_data(927) <= "010110111100";
rom_data(928) <= "010110111101";
rom_data(929) <= "010110111101";
rom_data(930) <= "010110111101";
rom_data(931) <= "010110111110";
rom_data(932) <= "010110111110";
rom_data(933) <= "010110111111";
rom_data(934) <= "010110111111";
rom_data(935) <= "010110111111";
rom_data(936) <= "010111000000";
rom_data(937) <= "010111000000";
rom_data(938) <= "010111000000";
rom_data(939) <= "010111000001";
rom_data(940) <= "010111000001";
rom_data(941) <= "010111000001";
rom_data(942) <= "010111000010";
rom_data(943) <= "010111000010";
rom_data(944) <= "010111000011";
rom_data(945) <= "010111000011";
rom_data(946) <= "010111000011";
rom_data(947) <= "010111000100";
rom_data(948) <= "010111000100";
rom_data(949) <= "010111000100";
rom_data(950) <= "010111000101";
rom_data(951) <= "010111000101";
rom_data(952) <= "010111000101";
rom_data(953) <= "010111000110";
rom_data(954) <= "010111000110";
rom_data(955) <= "010111000111";
rom_data(956) <= "010111000111";
rom_data(957) <= "010111000111";
rom_data(958) <= "010111001000";
rom_data(959) <= "010111001000";
rom_data(960) <= "010111001000";
rom_data(961) <= "010111001001";
rom_data(962) <= "010111001001";
rom_data(963) <= "010111001001";
rom_data(964) <= "010111001010";
rom_data(965) <= "010111001010";
rom_data(966) <= "010111001011";
rom_data(967) <= "010111001011";
rom_data(968) <= "010111001011";
rom_data(969) <= "010111001100";
rom_data(970) <= "010111001100";
rom_data(971) <= "010111001100";
rom_data(972) <= "010111001101";
rom_data(973) <= "010111001101";
rom_data(974) <= "010111001110";
rom_data(975) <= "010111001110";
rom_data(976) <= "010111001110";
rom_data(977) <= "010111001111";
rom_data(978) <= "010111001111";
rom_data(979) <= "010111001111";
rom_data(980) <= "010111010000";
rom_data(981) <= "010111010000";
rom_data(982) <= "010111010001";
rom_data(983) <= "010111010001";
rom_data(984) <= "010111010001";
rom_data(985) <= "010111010010";
rom_data(986) <= "010111010010";
rom_data(987) <= "010111010011";
rom_data(988) <= "010111010011";
rom_data(989) <= "010111010011";
rom_data(990) <= "010111010100";
rom_data(991) <= "010111010100";
rom_data(992) <= "010111010100";
rom_data(993) <= "010111010101";
rom_data(994) <= "010111010101";
rom_data(995) <= "010111010110";
rom_data(996) <= "010111010110";
rom_data(997) <= "010111010110";
rom_data(998) <= "010111010111";
rom_data(999) <= "010111010111";
rom_data(1000) <= "010111011000";
rom_data(1001) <= "010111011000";
rom_data(1002) <= "010111011000";
rom_data(1003) <= "010111011001";
rom_data(1004) <= "010111011001";
rom_data(1005) <= "010111011001";
rom_data(1006) <= "010111011010";
rom_data(1007) <= "010111011010";
rom_data(1008) <= "010111011011";
rom_data(1009) <= "010111011011";
rom_data(1010) <= "010111011011";
rom_data(1011) <= "010111011100";
rom_data(1012) <= "010111011100";
rom_data(1013) <= "010111011101";
rom_data(1014) <= "010111011101";
rom_data(1015) <= "010111011101";
rom_data(1016) <= "010111011110";
rom_data(1017) <= "010111011110";
rom_data(1018) <= "010111011111";
rom_data(1019) <= "010111011111";
rom_data(1020) <= "010111011111";
rom_data(1021) <= "010111100000";
rom_data(1022) <= "010111100000";
rom_data(1023) <= "010111100001";


process(i_clk)
begin
	if rising_edge(i_clk) then
		if conv_integer(i_addr) < 1024 then
			o_data <= rom_data(conv_integer(i_addr));
		else
			o_data <= (others => '0');
		end if;
	end if;
end process;



end Behavioral;


